magic
tech scmos
magscale 1 2
timestamp 1736168001
<< metal1 >>
rect 298 814 310 816
rect 283 806 285 814
rect 293 806 295 814
rect 303 806 305 814
rect 313 806 315 814
rect 323 806 325 814
rect 298 804 310 806
rect 269 697 444 703
rect 509 677 579 683
rect 1069 677 1100 683
rect 413 657 428 663
rect 500 657 515 663
rect 212 637 254 643
rect 573 637 588 643
rect 1012 636 1016 644
rect 778 614 790 616
rect 763 606 765 614
rect 773 606 775 614
rect 783 606 785 614
rect 793 606 795 614
rect 803 606 805 614
rect 778 604 790 606
rect 532 557 563 563
rect 188 543 196 548
rect 188 537 211 543
rect 900 537 915 543
rect 116 517 131 523
rect 477 517 515 523
rect 525 517 588 523
rect 477 504 483 517
rect 788 517 899 523
rect 349 497 387 503
rect 298 414 310 416
rect 283 406 285 414
rect 293 406 295 414
rect 303 406 305 414
rect 313 406 315 414
rect 323 406 325 414
rect 298 404 310 406
rect 749 377 812 383
rect 1066 376 1068 384
rect 772 357 835 363
rect 148 337 163 343
rect 412 332 420 336
rect 125 317 140 323
rect 413 317 451 323
rect 84 297 99 303
rect 605 297 652 303
rect 109 277 131 283
rect 468 277 483 283
rect 621 277 636 283
rect 778 214 790 216
rect 763 206 765 214
rect 773 206 775 214
rect 783 206 785 214
rect 793 206 795 214
rect 803 206 805 214
rect 778 204 790 206
rect 1069 177 1084 183
rect 317 157 387 163
rect 317 143 323 157
rect 548 156 556 164
rect 301 137 323 143
rect 472 136 476 144
rect 573 137 611 143
rect 589 117 604 123
rect 637 117 675 123
rect 669 104 675 117
rect 988 117 1011 123
rect 988 114 996 117
rect 404 97 419 103
rect 429 97 444 103
rect 708 97 723 103
rect 298 14 310 16
rect 283 6 285 14
rect 293 6 295 14
rect 303 6 305 14
rect 313 6 315 14
rect 323 6 325 14
rect 298 4 310 6
<< m2contact >>
rect 275 806 283 814
rect 285 806 293 814
rect 295 806 303 814
rect 305 806 313 814
rect 315 806 323 814
rect 325 806 333 814
rect 76 696 84 704
rect 444 696 452 704
rect 492 696 500 704
rect 652 696 660 704
rect 844 696 852 704
rect 284 676 292 684
rect 668 676 676 684
rect 796 676 804 684
rect 972 676 980 684
rect 1100 676 1108 684
rect 60 656 68 664
rect 300 656 308 664
rect 428 656 436 664
rect 492 656 500 664
rect 524 656 532 664
rect 556 656 564 664
rect 668 656 676 664
rect 828 656 836 664
rect 188 636 196 644
rect 204 636 212 644
rect 508 636 516 644
rect 588 636 596 644
rect 636 636 644 644
rect 956 636 964 644
rect 1004 636 1012 644
rect 755 606 763 614
rect 765 606 773 614
rect 775 606 783 614
rect 785 606 793 614
rect 795 606 803 614
rect 805 606 813 614
rect 188 576 196 584
rect 380 576 388 584
rect 60 556 68 564
rect 492 556 500 564
rect 524 556 532 564
rect 732 556 740 564
rect 860 556 868 564
rect 940 556 948 564
rect 364 536 372 544
rect 412 536 420 544
rect 428 536 436 544
rect 460 536 468 544
rect 572 536 580 544
rect 604 536 612 544
rect 668 536 676 544
rect 764 536 772 544
rect 892 536 900 544
rect 972 536 980 544
rect 1004 536 1012 544
rect 76 516 84 524
rect 108 516 116 524
rect 220 516 228 524
rect 236 516 244 524
rect 444 516 452 524
rect 588 516 596 524
rect 684 516 692 524
rect 700 516 708 524
rect 748 516 756 524
rect 780 516 788 524
rect 956 516 964 524
rect 1020 516 1028 524
rect 1052 516 1060 524
rect 252 496 260 504
rect 332 496 340 504
rect 476 496 484 504
rect 716 496 724 504
rect 1036 496 1044 504
rect 1068 476 1076 484
rect 1004 456 1012 464
rect 1052 456 1060 464
rect 940 436 948 444
rect 275 406 283 414
rect 285 406 293 414
rect 295 406 303 414
rect 305 406 313 414
rect 315 406 323 414
rect 325 406 333 414
rect 44 376 52 384
rect 220 376 228 384
rect 476 376 484 384
rect 540 376 548 384
rect 812 376 820 384
rect 1020 376 1028 384
rect 1068 376 1076 384
rect 764 356 772 364
rect 28 336 36 344
rect 140 336 148 344
rect 172 336 180 344
rect 412 336 420 344
rect 524 336 532 344
rect 732 336 740 344
rect 956 336 964 344
rect 60 316 68 324
rect 76 316 84 324
rect 140 316 148 324
rect 204 316 212 324
rect 460 316 468 324
rect 556 316 564 324
rect 572 316 580 324
rect 684 316 692 324
rect 700 316 708 324
rect 908 316 916 324
rect 924 316 932 324
rect 972 316 980 324
rect 1036 316 1044 324
rect 44 296 52 304
rect 76 296 84 304
rect 188 296 196 304
rect 252 296 260 304
rect 540 296 548 304
rect 652 296 660 304
rect 716 296 724 304
rect 876 296 884 304
rect 940 296 948 304
rect 988 296 996 304
rect 1068 296 1076 304
rect 268 276 276 284
rect 380 276 388 284
rect 460 276 468 284
rect 492 276 500 284
rect 572 276 580 284
rect 636 276 644 284
rect 684 276 692 284
rect 860 276 868 284
rect 908 276 916 284
rect 1084 276 1092 284
rect 140 256 148 264
rect 236 256 244 264
rect 300 256 308 264
rect 428 256 436 264
rect 844 256 852 264
rect 284 236 292 244
rect 412 236 420 244
rect 755 206 763 214
rect 765 206 773 214
rect 775 206 783 214
rect 785 206 793 214
rect 795 206 803 214
rect 805 206 813 214
rect 988 176 996 184
rect 1084 176 1092 184
rect 108 156 116 164
rect 396 156 404 164
rect 540 156 548 164
rect 732 156 740 164
rect 860 156 868 164
rect 1052 156 1060 164
rect 444 136 452 144
rect 476 136 484 144
rect 540 136 548 144
rect 652 136 660 144
rect 700 136 708 144
rect 44 116 52 124
rect 124 116 132 124
rect 268 116 276 124
rect 284 116 292 124
rect 492 116 500 124
rect 524 116 532 124
rect 604 116 612 124
rect 684 116 692 124
rect 876 116 884 124
rect 252 96 260 104
rect 396 96 404 104
rect 444 96 452 104
rect 508 96 516 104
rect 604 96 612 104
rect 668 96 676 104
rect 700 96 708 104
rect 12 76 20 84
rect 236 76 244 84
rect 476 76 484 84
rect 1036 36 1044 44
rect 275 6 283 14
rect 285 6 293 14
rect 295 6 303 14
rect 305 6 313 14
rect 315 6 323 14
rect 325 6 333 14
<< metal2 >>
rect 298 814 310 816
rect 283 806 285 814
rect 293 806 295 814
rect 303 806 305 814
rect 313 806 315 814
rect 323 806 325 814
rect 298 804 310 806
rect 61 644 67 656
rect 189 644 195 656
rect 61 564 67 636
rect 61 524 67 556
rect 77 444 83 516
rect 45 384 51 436
rect 29 344 35 376
rect 61 324 67 336
rect 77 324 83 396
rect 109 164 115 516
rect 173 344 179 516
rect 205 464 211 636
rect 381 584 387 696
rect 525 664 531 676
rect 429 584 435 656
rect 413 544 419 556
rect 429 544 435 576
rect 493 564 499 656
rect 509 584 515 636
rect 461 544 467 556
rect 221 504 227 516
rect 205 404 211 456
rect 221 384 227 496
rect 237 384 243 516
rect 253 504 259 536
rect 349 504 355 536
rect 365 524 371 536
rect 298 414 310 416
rect 283 406 285 414
rect 293 406 295 414
rect 303 406 305 414
rect 313 406 315 414
rect 323 406 325 414
rect 298 404 310 406
rect 205 324 211 356
rect 413 344 419 356
rect 253 304 259 316
rect 269 284 275 336
rect 141 264 147 276
rect 301 264 307 336
rect 445 324 451 516
rect 477 384 483 476
rect 509 344 515 576
rect 525 564 531 656
rect 589 524 595 636
rect 637 564 643 636
rect 525 344 531 456
rect 541 384 547 436
rect 461 304 467 316
rect 381 284 387 296
rect 237 244 243 256
rect 45 104 51 116
rect 253 104 259 156
rect 285 124 291 236
rect 397 104 403 156
rect 13 84 19 96
rect 237 84 243 96
rect 413 84 419 236
rect 445 144 451 296
rect 493 284 499 316
rect 493 264 499 276
rect 493 124 499 236
rect 525 124 531 336
rect 605 324 611 536
rect 580 317 595 323
rect 557 304 563 316
rect 541 284 547 296
rect 589 144 595 317
rect 605 124 611 316
rect 637 284 643 396
rect 653 364 659 696
rect 669 684 675 863
rect 1005 824 1011 863
rect 669 544 675 656
rect 797 644 803 676
rect 778 614 790 616
rect 763 606 765 614
rect 773 606 775 614
rect 783 606 785 614
rect 793 606 795 614
rect 803 606 805 614
rect 778 604 790 606
rect 685 524 691 536
rect 733 484 739 556
rect 781 504 787 516
rect 813 384 819 496
rect 653 304 659 356
rect 733 324 739 336
rect 685 304 691 316
rect 717 284 723 296
rect 733 164 739 296
rect 778 214 790 216
rect 763 206 765 214
rect 773 206 775 214
rect 783 206 785 214
rect 793 206 795 214
rect 803 206 805 214
rect 778 204 790 206
rect 829 164 835 656
rect 845 384 851 696
rect 861 564 867 676
rect 973 624 979 676
rect 861 404 867 556
rect 893 544 899 556
rect 893 524 899 536
rect 861 284 867 396
rect 909 324 915 616
rect 941 564 947 576
rect 1005 563 1011 636
rect 989 557 1011 563
rect 941 484 947 556
rect 957 524 963 556
rect 941 344 947 436
rect 989 364 995 557
rect 1005 484 1011 536
rect 1053 504 1059 516
rect 1021 423 1027 476
rect 1037 444 1043 496
rect 1053 464 1059 476
rect 1069 464 1075 476
rect 1005 417 1027 423
rect 957 344 963 356
rect 925 324 931 336
rect 957 324 963 336
rect 909 304 915 316
rect 877 264 883 296
rect 941 284 947 296
rect 845 204 851 256
rect 298 14 310 16
rect 283 6 285 14
rect 293 6 295 14
rect 303 6 305 14
rect 313 6 315 14
rect 323 6 325 14
rect 298 4 310 6
rect 973 -23 979 296
rect 989 184 995 196
rect 1005 124 1011 417
rect 1021 384 1027 396
rect 1053 304 1059 416
rect 1069 304 1075 336
rect 1053 164 1059 296
rect 1085 264 1091 276
rect 1085 184 1091 256
rect 1101 144 1107 676
rect 1037 -17 1043 36
rect 1021 -23 1043 -17
<< m3contact >>
rect 275 806 283 814
rect 285 806 293 814
rect 295 806 303 814
rect 305 806 313 814
rect 315 806 323 814
rect 325 806 333 814
rect 76 696 84 704
rect 380 696 388 704
rect 444 696 452 704
rect 492 696 500 704
rect 284 676 292 684
rect 188 656 196 664
rect 300 656 308 664
rect 60 636 68 644
rect 188 576 196 584
rect 60 516 68 524
rect 172 516 180 524
rect 44 436 52 444
rect 76 436 84 444
rect 76 396 84 404
rect 28 376 36 384
rect 60 336 68 344
rect 44 296 52 304
rect 76 296 84 304
rect 524 676 532 684
rect 556 656 564 664
rect 428 576 436 584
rect 412 556 420 564
rect 508 576 516 584
rect 460 556 468 564
rect 252 536 260 544
rect 348 536 356 544
rect 428 536 436 544
rect 220 496 228 504
rect 204 456 212 464
rect 204 396 212 404
rect 364 516 372 524
rect 332 496 340 504
rect 348 496 356 504
rect 275 406 283 414
rect 285 406 293 414
rect 295 406 303 414
rect 305 406 313 414
rect 315 406 323 414
rect 325 406 333 414
rect 236 376 244 384
rect 204 356 212 364
rect 412 356 420 364
rect 140 336 148 344
rect 172 336 180 344
rect 268 336 276 344
rect 300 336 308 344
rect 140 316 148 324
rect 252 316 260 324
rect 188 296 196 304
rect 140 276 148 284
rect 476 496 484 504
rect 476 476 484 484
rect 572 536 580 544
rect 636 556 644 564
rect 524 456 532 464
rect 540 436 548 444
rect 508 336 516 344
rect 524 336 532 344
rect 444 316 452 324
rect 492 316 500 324
rect 380 296 388 304
rect 444 296 452 304
rect 460 296 468 304
rect 428 256 436 264
rect 236 236 244 244
rect 252 156 260 164
rect 124 116 132 124
rect 268 116 276 124
rect 12 96 20 104
rect 44 96 52 104
rect 236 96 244 104
rect 396 96 404 104
rect 460 276 468 284
rect 492 256 500 264
rect 492 236 500 244
rect 476 136 484 144
rect 636 396 644 404
rect 572 316 580 324
rect 556 296 564 304
rect 540 276 548 284
rect 572 276 580 284
rect 540 156 548 164
rect 604 316 612 324
rect 540 136 548 144
rect 588 136 596 144
rect 1004 816 1012 824
rect 668 676 676 684
rect 668 656 676 664
rect 796 636 804 644
rect 755 606 763 614
rect 765 606 773 614
rect 775 606 783 614
rect 785 606 793 614
rect 795 606 803 614
rect 805 606 813 614
rect 684 536 692 544
rect 700 516 708 524
rect 716 496 724 504
rect 764 536 772 544
rect 748 516 756 524
rect 780 496 788 504
rect 812 496 820 504
rect 732 476 740 484
rect 652 356 660 364
rect 764 356 772 364
rect 700 316 708 324
rect 732 316 740 324
rect 684 296 692 304
rect 732 296 740 304
rect 684 276 692 284
rect 716 276 724 284
rect 755 206 763 214
rect 765 206 773 214
rect 775 206 783 214
rect 785 206 793 214
rect 795 206 803 214
rect 805 206 813 214
rect 860 676 868 684
rect 1100 676 1108 684
rect 956 636 964 644
rect 908 616 916 624
rect 972 616 980 624
rect 892 556 900 564
rect 892 516 900 524
rect 860 396 868 404
rect 844 376 852 384
rect 940 576 948 584
rect 956 556 964 564
rect 972 536 980 544
rect 940 476 948 484
rect 1020 516 1028 524
rect 1052 496 1060 504
rect 1004 476 1012 484
rect 1020 476 1028 484
rect 1004 456 1012 464
rect 1052 476 1060 484
rect 1068 456 1076 464
rect 1036 436 1044 444
rect 956 356 964 364
rect 988 356 996 364
rect 924 336 932 344
rect 940 336 948 344
rect 956 316 964 324
rect 972 316 980 324
rect 908 296 916 304
rect 972 296 980 304
rect 988 296 996 304
rect 908 276 916 284
rect 940 276 948 284
rect 876 256 884 264
rect 844 196 852 204
rect 828 156 836 164
rect 860 156 868 164
rect 652 136 660 144
rect 700 136 708 144
rect 492 116 500 124
rect 684 116 692 124
rect 876 116 884 124
rect 444 96 452 104
rect 508 96 516 104
rect 604 96 612 104
rect 668 96 676 104
rect 700 96 708 104
rect 412 76 420 84
rect 476 76 484 84
rect 275 6 283 14
rect 285 6 293 14
rect 295 6 303 14
rect 305 6 313 14
rect 315 6 323 14
rect 325 6 333 14
rect 988 196 996 204
rect 1052 416 1060 424
rect 1020 396 1028 404
rect 1036 316 1044 324
rect 1068 376 1076 384
rect 1068 336 1076 344
rect 1052 296 1060 304
rect 1084 256 1092 264
rect 1100 136 1108 144
rect 1004 116 1012 124
<< metal3 >>
rect 1012 817 1036 823
rect 274 814 334 816
rect 274 806 275 814
rect 284 806 285 814
rect 323 806 324 814
rect 333 806 334 814
rect 274 804 334 806
rect 84 697 380 703
rect 452 697 492 703
rect 292 677 524 683
rect 532 677 668 683
rect 676 677 860 683
rect 1108 677 1139 683
rect 196 657 300 663
rect 308 657 556 663
rect 564 657 668 663
rect 68 637 796 643
rect 964 637 1004 643
rect 916 617 972 623
rect 754 614 814 616
rect 754 606 755 614
rect 764 606 765 614
rect 803 606 804 614
rect 813 606 814 614
rect 754 604 814 606
rect 196 577 428 583
rect 516 577 940 583
rect 420 557 460 563
rect 644 557 883 563
rect 260 537 348 543
rect 436 537 572 543
rect 580 537 684 543
rect 692 537 764 543
rect 877 543 883 557
rect 900 557 956 563
rect 877 537 972 543
rect -35 517 60 523
rect 180 517 364 523
rect 372 517 700 523
rect 756 517 892 523
rect 948 517 1020 523
rect 228 497 332 503
rect 356 497 476 503
rect 724 497 780 503
rect 820 497 1052 503
rect 484 477 732 483
rect 948 477 1004 483
rect 1028 477 1052 483
rect 212 457 524 463
rect 1012 457 1068 463
rect 52 437 76 443
rect 548 437 1036 443
rect 1012 417 1052 423
rect 274 414 334 416
rect 274 406 275 414
rect 284 406 285 414
rect 323 406 324 414
rect 333 406 334 414
rect 274 404 334 406
rect 84 397 204 403
rect 644 397 860 403
rect 1028 397 1036 403
rect 36 377 236 383
rect 852 377 1068 383
rect 212 357 412 363
rect 660 357 764 363
rect 964 357 988 363
rect 68 337 140 343
rect 180 337 268 343
rect 308 337 508 343
rect 532 337 924 343
rect 948 337 1068 343
rect 148 317 252 323
rect 260 317 444 323
rect 500 317 572 323
rect 612 317 700 323
rect 740 317 956 323
rect 980 317 1036 323
rect 52 297 76 303
rect 196 297 380 303
rect 388 297 444 303
rect 452 297 460 303
rect 468 297 556 303
rect 564 297 684 303
rect 692 297 732 303
rect 740 297 908 303
rect 916 297 972 303
rect 996 297 1052 303
rect 148 277 460 283
rect 548 277 572 283
rect 692 277 716 283
rect 916 277 940 283
rect 436 257 492 263
rect 884 257 1084 263
rect 244 237 492 243
rect 754 214 814 216
rect 754 206 755 214
rect 764 206 765 214
rect 803 206 804 214
rect 813 206 814 214
rect 754 204 814 206
rect 852 197 940 203
rect 948 197 988 203
rect 260 157 540 163
rect 836 157 860 163
rect 484 137 540 143
rect 596 137 652 143
rect 660 137 700 143
rect 708 137 1100 143
rect 132 117 268 123
rect 500 117 684 123
rect 884 117 1004 123
rect -35 97 12 103
rect 52 97 236 103
rect 244 97 396 103
rect 452 97 508 103
rect 516 97 604 103
rect 676 97 700 103
rect 420 77 476 83
rect 274 14 334 16
rect 274 6 275 14
rect 284 6 285 14
rect 323 6 324 14
rect 333 6 334 14
rect 274 4 334 6
<< m4contact >>
rect 1036 816 1044 824
rect 276 806 283 814
rect 283 806 284 814
rect 288 806 293 814
rect 293 806 295 814
rect 295 806 296 814
rect 300 806 303 814
rect 303 806 305 814
rect 305 806 308 814
rect 312 806 313 814
rect 313 806 315 814
rect 315 806 320 814
rect 324 806 325 814
rect 325 806 332 814
rect 1004 636 1012 644
rect 756 606 763 614
rect 763 606 764 614
rect 768 606 773 614
rect 773 606 775 614
rect 775 606 776 614
rect 780 606 783 614
rect 783 606 785 614
rect 785 606 788 614
rect 792 606 793 614
rect 793 606 795 614
rect 795 606 800 614
rect 804 606 805 614
rect 805 606 812 614
rect 940 516 948 524
rect 1004 416 1012 424
rect 276 406 283 414
rect 283 406 284 414
rect 288 406 293 414
rect 293 406 295 414
rect 295 406 296 414
rect 300 406 303 414
rect 303 406 305 414
rect 305 406 308 414
rect 312 406 313 414
rect 313 406 315 414
rect 315 406 320 414
rect 324 406 325 414
rect 325 406 332 414
rect 1036 396 1044 404
rect 756 206 763 214
rect 763 206 764 214
rect 768 206 773 214
rect 773 206 775 214
rect 775 206 776 214
rect 780 206 783 214
rect 783 206 785 214
rect 785 206 788 214
rect 792 206 793 214
rect 793 206 795 214
rect 795 206 800 214
rect 804 206 805 214
rect 805 206 812 214
rect 940 196 948 204
rect 276 6 283 14
rect 283 6 284 14
rect 288 6 293 14
rect 293 6 295 14
rect 295 6 296 14
rect 300 6 303 14
rect 303 6 305 14
rect 305 6 308 14
rect 312 6 313 14
rect 313 6 315 14
rect 315 6 320 14
rect 324 6 325 14
rect 325 6 332 14
<< metal4 >>
rect 1034 824 1046 826
rect 1034 816 1036 824
rect 1044 816 1046 824
rect 272 814 336 816
rect 272 806 276 814
rect 284 806 288 814
rect 296 806 300 814
rect 308 806 312 814
rect 320 806 324 814
rect 332 806 336 814
rect 272 414 336 806
rect 272 406 276 414
rect 284 406 288 414
rect 296 406 300 414
rect 308 406 312 414
rect 320 406 324 414
rect 332 406 336 414
rect 272 14 336 406
rect 272 6 276 14
rect 284 6 288 14
rect 296 6 300 14
rect 308 6 312 14
rect 320 6 324 14
rect 332 6 336 14
rect 272 -10 336 6
rect 752 614 816 816
rect 752 606 756 614
rect 764 606 768 614
rect 776 606 780 614
rect 788 606 792 614
rect 800 606 804 614
rect 812 606 816 614
rect 752 214 816 606
rect 1002 644 1014 646
rect 1002 636 1004 644
rect 1012 636 1014 644
rect 752 206 756 214
rect 764 206 768 214
rect 776 206 780 214
rect 788 206 792 214
rect 800 206 804 214
rect 812 206 816 214
rect 752 -10 816 206
rect 938 524 950 526
rect 938 516 940 524
rect 948 516 950 524
rect 938 204 950 516
rect 1002 424 1014 636
rect 1002 416 1004 424
rect 1012 416 1014 424
rect 1002 414 1014 416
rect 1034 404 1046 816
rect 1034 396 1036 404
rect 1044 396 1046 404
rect 1034 394 1046 396
rect 938 196 940 204
rect 948 196 950 204
rect 938 194 950 196
use INVX1  _44_
timestamp 0
transform -1 0 744 0 -1 210
box -4 -6 36 206
use NAND2X1  _45_
timestamp 0
transform -1 0 712 0 -1 210
box -4 -6 52 206
use INVX1  _46_
timestamp 0
transform -1 0 248 0 1 210
box -4 -6 36 206
use INVX1  _47_
timestamp 0
transform 1 0 856 0 -1 610
box -4 -6 36 206
use OAI21X1  _48_
timestamp 0
transform 1 0 664 0 -1 610
box -4 -6 68 206
use NAND2X1  _49_
timestamp 0
transform -1 0 376 0 -1 610
box -4 -6 52 206
use INVX1  _50_
timestamp 0
transform 1 0 552 0 1 610
box -4 -6 36 206
use NOR2X1  _51_
timestamp 0
transform 1 0 488 0 -1 610
box -4 -6 52 206
use NAND2X1  _52_
timestamp 0
transform -1 0 504 0 1 210
box -4 -6 52 206
use INVX1  _53_
timestamp 0
transform -1 0 152 0 1 210
box -4 -6 36 206
use OAI21X1  _54_
timestamp 0
transform 1 0 424 0 -1 610
box -4 -6 68 206
use NAND2X1  _55_
timestamp 0
transform -1 0 424 0 -1 610
box -4 -6 52 206
use INVX1  _56_
timestamp 0
transform -1 0 424 0 1 610
box -4 -6 36 206
use NOR3X1  _57_
timestamp 0
transform -1 0 328 0 1 610
box -4 -6 132 206
use NAND2X1  _58_
timestamp 0
transform -1 0 120 0 1 210
box -4 -6 52 206
use INVX1  _59_
timestamp 0
transform 1 0 424 0 1 210
box -4 -6 36 206
use NAND3X1  _60_
timestamp 0
transform -1 0 216 0 1 210
box -4 -6 68 206
use OAI21X1  _61_
timestamp 0
transform 1 0 200 0 -1 610
box -4 -6 68 206
use NAND3X1  _62_
timestamp 0
transform -1 0 72 0 1 210
box -4 -6 68 206
use INVX1  _63_
timestamp 0
transform -1 0 856 0 1 210
box -4 -6 36 206
use OAI21X1  _64_
timestamp 0
transform -1 0 632 0 1 210
box -4 -6 68 206
use NAND3X1  _65_
timestamp 0
transform -1 0 568 0 1 210
box -4 -6 68 206
use NOR3X1  _66_
timestamp 0
transform 1 0 536 0 -1 610
box -4 -6 132 206
use XNOR2X1  _67_
timestamp 0
transform -1 0 1080 0 1 610
box -4 -6 116 206
use OAI21X1  _68_
timestamp 0
transform 1 0 632 0 1 210
box -4 -6 68 206
use NAND3X1  _69_
timestamp 0
transform 1 0 696 0 1 210
box -4 -6 68 206
use NOR3X1  _70_
timestamp 0
transform -1 0 552 0 1 610
box -4 -6 132 206
use AOI21X1  _71_
timestamp 0
transform -1 0 792 0 -1 610
box -4 -6 68 206
use NOR3X1  _72_
timestamp 0
transform -1 0 712 0 1 610
box -4 -6 132 206
use AOI22X1  _73_
timestamp 0
transform 1 0 952 0 -1 610
box -4 -6 84 206
use NAND3X1  _74_
timestamp 0
transform 1 0 1032 0 -1 610
box -4 -6 68 206
use INVX1  _75_
timestamp 0
transform 1 0 1048 0 -1 210
box -4 -6 36 206
use OAI21X1  _76_
timestamp 0
transform 1 0 856 0 1 210
box -4 -6 68 206
use NAND3X1  _77_
timestamp 0
transform 1 0 920 0 1 210
box -4 -6 68 206
use AOI21X1  _78_
timestamp 0
transform 1 0 888 0 -1 610
box -4 -6 68 206
use OAI21X1  _79_
timestamp 0
transform -1 0 1096 0 1 210
box -4 -6 68 206
use INVX1  _80_
timestamp 0
transform -1 0 408 0 -1 210
box -4 -6 36 206
use AOI21X1  _81_
timestamp 0
transform 1 0 248 0 1 210
box -4 -6 68 206
use NAND2X1  _82_
timestamp 0
transform -1 0 456 0 -1 210
box -4 -6 52 206
use OAI21X1  _83_
timestamp 0
transform -1 0 664 0 -1 210
box -4 -6 68 206
use NAND2X1  _84_
timestamp 0
transform 1 0 376 0 1 210
box -4 -6 52 206
use NAND3X1  _85_
timestamp 0
transform -1 0 520 0 -1 210
box -4 -6 68 206
use AOI22X1  _86_
timestamp 0
transform -1 0 600 0 -1 210
box -4 -6 84 206
use OAI21X1  _87_
timestamp 0
transform -1 0 312 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _88_
timestamp 0
transform 1 0 8 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _89_
timestamp 0
transform 1 0 56 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _90_
timestamp 0
transform 1 0 808 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _91_
timestamp 0
transform 1 0 776 0 1 610
box -4 -6 196 206
use DFFPOSX1  _92_
timestamp 0
transform 1 0 8 0 1 610
box -4 -6 196 206
use BUFX2  _93_
timestamp 0
transform 1 0 1000 0 -1 210
box -4 -6 52 206
use BUFX2  _94_
timestamp 0
transform 1 0 984 0 1 210
box -4 -6 52 206
use BUFX2  _95_
timestamp 0
transform -1 0 56 0 -1 210
box -4 -6 52 206
use FILL  FILL9520x100
timestamp 0
transform -1 0 1096 0 -1 210
box -4 -6 20 206
use FILL  FILL9520x6100
timestamp 0
transform 1 0 1080 0 1 610
box -4 -6 20 206
use FILL  SFILL2640x4100
timestamp 0
transform -1 0 280 0 -1 610
box -4 -6 20 206
use FILL  SFILL2800x4100
timestamp 0
transform -1 0 296 0 -1 610
box -4 -6 20 206
use FILL  SFILL2960x4100
timestamp 0
transform -1 0 312 0 -1 610
box -4 -6 20 206
use FILL  SFILL3120x100
timestamp 0
transform -1 0 328 0 -1 210
box -4 -6 20 206
use FILL  SFILL3120x2100
timestamp 0
transform 1 0 312 0 1 210
box -4 -6 20 206
use FILL  SFILL3120x4100
timestamp 0
transform -1 0 328 0 -1 610
box -4 -6 20 206
use FILL  SFILL3280x100
timestamp 0
transform -1 0 344 0 -1 210
box -4 -6 20 206
use FILL  SFILL3280x2100
timestamp 0
transform 1 0 328 0 1 210
box -4 -6 20 206
use FILL  SFILL3280x6100
timestamp 0
transform 1 0 328 0 1 610
box -4 -6 20 206
use FILL  SFILL3440x100
timestamp 0
transform -1 0 360 0 -1 210
box -4 -6 20 206
use FILL  SFILL3440x2100
timestamp 0
transform 1 0 344 0 1 210
box -4 -6 20 206
use FILL  SFILL3440x6100
timestamp 0
transform 1 0 344 0 1 610
box -4 -6 20 206
use FILL  SFILL3600x100
timestamp 0
transform -1 0 376 0 -1 210
box -4 -6 20 206
use FILL  SFILL3600x2100
timestamp 0
transform 1 0 360 0 1 210
box -4 -6 20 206
use FILL  SFILL3600x6100
timestamp 0
transform 1 0 360 0 1 610
box -4 -6 20 206
use FILL  SFILL3760x6100
timestamp 0
transform 1 0 376 0 1 610
box -4 -6 20 206
use FILL  SFILL7120x6100
timestamp 0
transform 1 0 712 0 1 610
box -4 -6 20 206
use FILL  SFILL7280x6100
timestamp 0
transform 1 0 728 0 1 610
box -4 -6 20 206
use FILL  SFILL7440x100
timestamp 0
transform -1 0 760 0 -1 210
box -4 -6 20 206
use FILL  SFILL7440x6100
timestamp 0
transform 1 0 744 0 1 610
box -4 -6 20 206
use FILL  SFILL7600x100
timestamp 0
transform -1 0 776 0 -1 210
box -4 -6 20 206
use FILL  SFILL7600x2100
timestamp 0
transform 1 0 760 0 1 210
box -4 -6 20 206
use FILL  SFILL7600x6100
timestamp 0
transform 1 0 760 0 1 610
box -4 -6 20 206
use FILL  SFILL7760x100
timestamp 0
transform -1 0 792 0 -1 210
box -4 -6 20 206
use FILL  SFILL7760x2100
timestamp 0
transform 1 0 776 0 1 210
box -4 -6 20 206
use FILL  SFILL7920x100
timestamp 0
transform -1 0 808 0 -1 210
box -4 -6 20 206
use FILL  SFILL7920x2100
timestamp 0
transform 1 0 792 0 1 210
box -4 -6 20 206
use FILL  SFILL7920x4100
timestamp 0
transform -1 0 808 0 -1 610
box -4 -6 20 206
use FILL  SFILL8080x2100
timestamp 0
transform 1 0 808 0 1 210
box -4 -6 20 206
use FILL  SFILL8080x4100
timestamp 0
transform -1 0 824 0 -1 610
box -4 -6 20 206
use FILL  SFILL8240x4100
timestamp 0
transform -1 0 840 0 -1 610
box -4 -6 20 206
use FILL  SFILL8400x4100
timestamp 0
transform -1 0 856 0 -1 610
box -4 -6 20 206
<< labels >>
flabel metal4 s 752 -10 816 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 272 -10 336 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 1005 857 1011 863 3 FreeSans 24 90 0 0 change[1]
port 2 nsew
flabel metal2 s 1021 -23 1027 -17 7 FreeSans 24 270 0 0 change[0]
port 3 nsew
flabel metal3 s -35 517 -29 523 7 FreeSans 24 0 0 0 clk
port 4 nsew
flabel metal2 s 973 -23 979 -17 7 FreeSans 24 270 0 0 in[1]
port 5 nsew
flabel metal3 s 1133 677 1139 683 3 FreeSans 24 0 0 0 in[0]
port 6 nsew
flabel metal3 s -35 97 -29 103 7 FreeSans 24 0 0 0 out
port 7 nsew
flabel metal2 s 669 857 675 863 3 FreeSans 24 90 0 0 rst
port 8 nsew
<< properties >>
string FIXED_BBOX -48 -40 1152 860
<< end >>
