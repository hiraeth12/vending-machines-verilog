VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vending_machine_18105070
  CLASS BLOCK ;
  FOREIGN vending_machine_18105070 ;
  ORIGIN 4.800 4.000 ;
  SIZE 120.000 BY 90.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 8.200 61.600 9.200 64.200 ;
        RECT 11.600 61.600 12.400 64.200 ;
        RECT 17.200 61.600 18.000 66.000 ;
        RECT 26.800 61.600 27.600 63.800 ;
        RECT 30.000 61.600 30.800 64.200 ;
        RECT 41.200 61.600 42.000 64.200 ;
        RECT 49.200 61.600 50.000 63.800 ;
        RECT 52.400 61.600 53.200 64.200 ;
        RECT 55.600 61.600 56.400 64.200 ;
        RECT 65.200 61.600 66.000 63.800 ;
        RECT 68.400 61.600 69.200 64.200 ;
        RECT 79.600 61.600 80.400 66.200 ;
        RECT 85.000 61.600 86.000 64.200 ;
        RECT 88.400 61.600 89.200 64.200 ;
        RECT 94.000 61.600 94.800 66.000 ;
        RECT 98.800 61.600 99.800 65.600 ;
        RECT 105.000 62.200 106.000 65.600 ;
        RECT 105.000 61.600 105.800 62.200 ;
        RECT 0.400 60.400 110.000 61.600 ;
        RECT 2.800 55.800 3.600 60.400 ;
        RECT 8.200 57.800 9.200 60.400 ;
        RECT 11.600 57.800 12.400 60.400 ;
        RECT 17.200 56.000 18.000 60.400 ;
        RECT 22.000 56.600 22.800 60.400 ;
        RECT 36.400 55.800 37.200 60.400 ;
        RECT 41.200 55.800 42.000 60.400 ;
        RECT 44.400 56.600 45.200 60.400 ;
        RECT 49.200 57.800 50.000 60.400 ;
        RECT 52.400 57.800 53.200 60.400 ;
        RECT 55.600 57.800 56.400 60.400 ;
        RECT 58.800 58.200 59.600 60.400 ;
        RECT 68.400 56.600 69.200 60.400 ;
        RECT 73.200 57.800 74.000 60.400 ;
        RECT 77.400 55.800 78.200 60.400 ;
        RECT 86.000 57.800 86.800 60.400 ;
        RECT 89.800 55.800 90.600 60.400 ;
        RECT 94.000 57.800 94.800 60.400 ;
        RECT 96.000 55.800 96.800 60.400 ;
        RECT 102.000 55.800 102.800 60.400 ;
        RECT 103.600 53.800 104.400 60.400 ;
        RECT 6.000 21.600 6.800 28.200 ;
        RECT 10.800 21.600 11.600 26.200 ;
        RECT 14.000 21.600 14.800 24.200 ;
        RECT 20.400 21.600 21.200 28.200 ;
        RECT 23.600 21.600 24.400 24.200 ;
        RECT 25.800 21.600 26.600 26.200 ;
        RECT 30.000 21.600 30.800 24.200 ;
        RECT 38.000 21.600 38.800 26.200 ;
        RECT 42.800 21.600 43.600 24.200 ;
        RECT 49.200 21.600 50.000 26.200 ;
        RECT 55.600 21.600 56.400 28.200 ;
        RECT 60.400 21.600 61.200 25.400 ;
        RECT 65.200 21.600 66.000 25.400 ;
        RECT 70.000 21.600 70.800 28.200 ;
        RECT 84.400 21.600 85.200 24.200 ;
        RECT 87.600 21.600 88.400 25.400 ;
        RECT 92.400 21.600 93.200 28.200 ;
        RECT 100.400 21.600 101.200 26.200 ;
        RECT 106.800 21.600 107.600 25.400 ;
        RECT 0.400 20.400 110.000 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 13.000 17.800 14.000 20.400 ;
        RECT 16.400 17.800 17.200 20.400 ;
        RECT 22.000 16.000 22.800 20.400 ;
        RECT 28.400 16.600 29.200 20.400 ;
        RECT 39.600 17.800 40.400 20.400 ;
        RECT 44.400 15.800 45.200 20.400 ;
        RECT 50.800 13.800 51.600 20.400 ;
        RECT 52.400 15.800 53.200 20.400 ;
        RECT 58.400 15.800 59.200 20.400 ;
        RECT 63.600 16.600 64.400 20.400 ;
        RECT 70.000 15.800 70.800 20.400 ;
        RECT 73.200 17.800 74.000 20.400 ;
        RECT 82.800 15.800 83.600 20.400 ;
        RECT 88.200 17.800 89.200 20.400 ;
        RECT 91.600 17.800 92.400 20.400 ;
        RECT 97.200 16.000 98.000 20.400 ;
        RECT 102.000 15.800 102.800 20.400 ;
        RECT 105.200 17.800 106.000 20.400 ;
      LAYER metal2 ;
        RECT 77.800 61.400 79.000 61.600 ;
        RECT 75.500 60.600 81.300 61.400 ;
        RECT 77.800 60.400 79.000 60.600 ;
        RECT 77.800 21.400 79.000 21.600 ;
        RECT 75.500 20.600 81.300 21.400 ;
        RECT 77.800 20.400 79.000 20.600 ;
      LAYER metal3 ;
        RECT 75.400 60.400 81.400 61.600 ;
        RECT 75.400 20.400 81.400 21.600 ;
      LAYER metal4 ;
        RECT 75.200 -1.000 81.600 81.600 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 80.400 110.000 81.600 ;
        RECT 2.800 72.000 3.600 80.400 ;
        RECT 8.400 75.800 9.200 80.400 ;
        RECT 11.600 75.800 12.400 80.400 ;
        RECT 17.200 71.800 18.000 80.400 ;
        RECT 30.000 73.800 30.800 80.400 ;
        RECT 41.200 75.800 42.000 80.400 ;
        RECT 52.400 73.800 53.200 80.400 ;
        RECT 55.600 75.800 56.400 80.400 ;
        RECT 68.400 73.800 69.200 80.400 ;
        RECT 79.600 72.000 80.400 80.400 ;
        RECT 85.200 75.800 86.000 80.400 ;
        RECT 88.400 75.800 89.200 80.400 ;
        RECT 94.000 71.800 94.800 80.400 ;
        RECT 98.800 73.200 99.800 80.400 ;
        RECT 105.000 79.800 105.800 80.400 ;
        RECT 105.000 73.200 106.000 79.800 ;
        RECT 2.800 41.600 3.600 50.000 ;
        RECT 8.400 41.600 9.200 46.200 ;
        RECT 11.600 41.600 12.400 46.200 ;
        RECT 17.200 41.600 18.000 50.200 ;
        RECT 20.400 41.600 21.200 50.200 ;
        RECT 24.600 41.600 25.400 46.200 ;
        RECT 33.200 41.600 34.000 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 38.000 41.600 38.800 46.200 ;
        RECT 41.200 41.600 42.000 46.200 ;
        RECT 42.800 41.600 43.600 50.200 ;
        RECT 47.000 41.600 47.800 46.200 ;
        RECT 49.200 41.600 50.000 50.200 ;
        RECT 55.600 41.600 56.400 48.200 ;
        RECT 66.800 41.600 67.600 50.200 ;
        RECT 71.000 41.600 71.800 46.200 ;
        RECT 76.400 41.600 77.200 49.000 ;
        RECT 86.000 41.600 86.800 46.200 ;
        RECT 90.800 41.600 91.600 49.000 ;
        RECT 97.200 41.600 98.000 49.000 ;
        RECT 103.600 41.600 104.400 46.200 ;
        RECT 106.800 41.600 107.600 45.800 ;
        RECT 0.400 40.400 110.000 41.600 ;
        RECT 2.800 36.200 3.600 40.400 ;
        RECT 6.000 35.800 6.800 40.400 ;
        RECT 7.600 35.800 8.400 40.400 ;
        RECT 10.800 35.800 11.600 40.400 ;
        RECT 14.000 35.800 14.800 40.400 ;
        RECT 17.200 36.200 18.000 40.400 ;
        RECT 20.400 35.800 21.200 40.400 ;
        RECT 23.600 35.800 24.400 40.400 ;
        RECT 26.800 33.000 27.600 40.400 ;
        RECT 38.000 35.800 38.800 40.400 ;
        RECT 41.200 35.800 42.000 40.400 ;
        RECT 42.800 35.800 43.600 40.400 ;
        RECT 46.000 35.800 46.800 40.400 ;
        RECT 49.200 35.800 50.000 40.400 ;
        RECT 52.400 36.200 53.200 40.400 ;
        RECT 55.600 35.800 56.400 40.400 ;
        RECT 57.800 35.800 58.600 40.400 ;
        RECT 62.000 31.800 62.800 40.400 ;
        RECT 63.600 31.800 64.400 40.400 ;
        RECT 67.800 35.800 68.600 40.400 ;
        RECT 70.000 35.800 70.800 40.400 ;
        RECT 73.200 36.200 74.000 40.400 ;
        RECT 84.400 35.800 85.200 40.400 ;
        RECT 86.000 31.800 86.800 40.400 ;
        RECT 90.200 35.800 91.000 40.400 ;
        RECT 92.400 35.800 93.200 40.400 ;
        RECT 95.600 36.200 96.400 40.400 ;
        RECT 100.400 33.000 101.200 40.400 ;
        RECT 104.200 35.800 105.000 40.400 ;
        RECT 108.400 31.800 109.200 40.400 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 7.600 1.600 8.400 10.000 ;
        RECT 13.200 1.600 14.000 6.200 ;
        RECT 16.400 1.600 17.200 6.200 ;
        RECT 22.000 1.600 22.800 10.200 ;
        RECT 25.800 1.600 26.600 6.200 ;
        RECT 30.000 1.600 30.800 10.200 ;
        RECT 39.600 1.600 40.400 6.200 ;
        RECT 41.200 1.600 42.000 6.200 ;
        RECT 44.400 1.600 45.200 6.200 ;
        RECT 47.600 1.600 48.400 5.800 ;
        RECT 50.800 1.600 51.600 6.200 ;
        RECT 57.200 1.600 58.000 9.000 ;
        RECT 61.000 1.600 61.800 6.200 ;
        RECT 65.200 1.600 66.000 10.200 ;
        RECT 66.800 1.600 67.600 6.200 ;
        RECT 70.000 1.600 70.800 6.200 ;
        RECT 73.200 1.600 74.000 6.200 ;
        RECT 82.800 1.600 83.600 10.000 ;
        RECT 88.400 1.600 89.200 6.200 ;
        RECT 91.600 1.600 92.400 6.200 ;
        RECT 97.200 1.600 98.000 10.200 ;
        RECT 102.000 1.600 102.800 9.000 ;
        RECT 105.200 1.600 106.000 6.200 ;
        RECT 0.400 0.400 110.000 1.600 ;
      LAYER metal2 ;
        RECT 29.800 81.400 31.000 81.600 ;
        RECT 27.500 80.600 33.300 81.400 ;
        RECT 29.800 80.400 31.000 80.600 ;
        RECT 29.800 41.400 31.000 41.600 ;
        RECT 27.500 40.600 33.300 41.400 ;
        RECT 29.800 40.400 31.000 40.600 ;
        RECT 29.800 1.400 31.000 1.600 ;
        RECT 27.500 0.600 33.300 1.400 ;
        RECT 29.800 0.400 31.000 0.600 ;
      LAYER metal3 ;
        RECT 27.400 80.400 33.400 81.600 ;
        RECT 27.400 40.400 33.400 41.600 ;
        RECT 27.400 0.400 33.400 1.600 ;
      LAYER metal4 ;
        RECT 27.200 -1.000 33.600 81.600 ;
    END
  END vdd
  PIN change[1]
    PORT
      LAYER metal1 ;
        RECT 102.000 31.800 102.800 39.800 ;
        RECT 102.200 29.600 102.800 31.800 ;
        RECT 102.000 22.200 102.800 29.600 ;
      LAYER metal2 ;
        RECT 100.500 82.400 101.100 86.300 ;
        RECT 100.400 81.600 101.200 82.400 ;
        RECT 102.000 39.600 102.800 40.400 ;
        RECT 102.100 38.400 102.700 39.600 ;
        RECT 102.000 37.600 102.800 38.400 ;
      LAYER metal3 ;
        RECT 100.400 82.300 101.200 82.400 ;
        RECT 103.600 82.300 104.400 82.400 ;
        RECT 100.400 81.700 104.400 82.300 ;
        RECT 100.400 81.600 101.200 81.700 ;
        RECT 103.600 81.600 104.400 81.700 ;
        RECT 102.000 40.300 102.800 40.400 ;
        RECT 103.600 40.300 104.400 40.400 ;
        RECT 102.000 39.700 104.400 40.300 ;
        RECT 102.000 39.600 102.800 39.700 ;
        RECT 103.600 39.600 104.400 39.700 ;
      LAYER metal4 ;
        RECT 103.400 39.400 104.600 82.600 ;
    END
  END change[1]
  PIN change[0]
    PORT
      LAYER metal1 ;
        RECT 103.600 12.400 104.400 19.800 ;
        RECT 103.800 10.200 104.400 12.400 ;
        RECT 103.600 2.200 104.400 10.200 ;
      LAYER metal2 ;
        RECT 103.600 3.600 104.400 4.400 ;
        RECT 103.700 -1.700 104.300 3.600 ;
        RECT 102.100 -2.300 104.300 -1.700 ;
    END
  END change[0]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 14.200 73.200 15.600 74.000 ;
        RECT 91.000 73.200 92.400 74.000 ;
        RECT 14.200 72.200 14.800 73.200 ;
        RECT 91.000 72.200 91.600 73.200 ;
        RECT 12.400 71.600 14.800 72.200 ;
        RECT 89.200 71.600 91.600 72.200 ;
        RECT 5.000 68.400 5.800 68.600 ;
        RECT 12.400 68.400 13.000 71.600 ;
        RECT 81.800 68.400 82.600 68.600 ;
        RECT 89.200 68.400 89.800 71.600 ;
        RECT 2.000 67.800 13.000 68.400 ;
        RECT 78.800 67.800 89.800 68.400 ;
        RECT 2.000 67.600 3.600 67.800 ;
        RECT 6.200 66.400 6.800 67.800 ;
        RECT 11.800 67.600 12.600 67.800 ;
        RECT 78.800 67.600 80.400 67.800 ;
        RECT 83.000 66.400 83.600 67.800 ;
        RECT 88.600 67.600 89.400 67.800 ;
        RECT 6.000 64.800 6.800 66.400 ;
        RECT 82.800 64.800 83.600 66.400 ;
        RECT 6.000 55.600 6.800 57.200 ;
        RECT 2.000 54.200 3.600 54.400 ;
        RECT 6.200 54.200 6.800 55.600 ;
        RECT 11.800 54.200 12.600 54.400 ;
        RECT 2.000 53.600 13.000 54.200 ;
        RECT 5.000 53.400 5.800 53.600 ;
        RECT 10.800 52.300 11.600 52.400 ;
        RECT 12.400 52.300 13.000 53.600 ;
        RECT 10.800 51.700 13.100 52.300 ;
        RECT 10.800 51.600 11.600 51.700 ;
        RECT 12.400 50.400 13.000 51.700 ;
        RECT 12.400 49.800 14.800 50.400 ;
        RECT 14.200 48.800 14.800 49.800 ;
        RECT 14.200 48.000 15.600 48.800 ;
        RECT 10.800 15.600 11.600 17.200 ;
        RECT 86.000 15.600 86.800 17.200 ;
        RECT 6.800 14.200 8.400 14.400 ;
        RECT 11.000 14.200 11.600 15.600 ;
        RECT 16.600 14.200 17.400 14.400 ;
        RECT 82.000 14.200 83.600 14.400 ;
        RECT 86.200 14.200 86.800 15.600 ;
        RECT 91.800 14.200 92.600 14.400 ;
        RECT 6.800 13.600 17.800 14.200 ;
        RECT 82.000 13.600 93.000 14.200 ;
        RECT 9.800 13.400 10.600 13.600 ;
        RECT 17.200 10.400 17.800 13.600 ;
        RECT 85.000 13.400 85.800 13.600 ;
        RECT 92.400 10.400 93.000 13.600 ;
        RECT 17.200 9.800 19.600 10.400 ;
        RECT 92.400 9.800 94.800 10.400 ;
        RECT 19.000 8.800 19.600 9.800 ;
        RECT 94.200 8.800 94.800 9.800 ;
        RECT 19.000 8.000 20.400 8.800 ;
        RECT 94.200 8.000 95.600 8.800 ;
      LAYER metal2 ;
        RECT 79.600 67.600 80.400 68.400 ;
        RECT 6.000 65.600 6.800 66.400 ;
        RECT 6.100 64.400 6.700 65.600 ;
        RECT 79.700 64.400 80.300 67.600 ;
        RECT 82.800 65.600 83.600 66.400 ;
        RECT 6.000 63.600 6.800 64.400 ;
        RECT 79.600 63.600 80.400 64.400 ;
        RECT 6.100 56.400 6.700 63.600 ;
        RECT 6.000 55.600 6.800 56.400 ;
        RECT 6.100 52.400 6.700 55.600 ;
        RECT 6.000 51.600 6.800 52.400 ;
        RECT 10.800 51.600 11.600 52.400 ;
        RECT 10.900 16.400 11.500 51.600 ;
        RECT 82.900 16.400 83.500 65.600 ;
        RECT 10.800 15.600 11.600 16.400 ;
        RECT 82.800 15.600 83.600 16.400 ;
        RECT 86.000 15.600 86.800 16.400 ;
      LAYER metal3 ;
        RECT 6.000 64.300 6.800 64.400 ;
        RECT 79.600 64.300 80.400 64.400 ;
        RECT 6.000 63.700 80.400 64.300 ;
        RECT 6.000 63.600 6.800 63.700 ;
        RECT 79.600 63.600 80.400 63.700 ;
        RECT 6.000 52.300 6.800 52.400 ;
        RECT -3.500 51.700 6.800 52.300 ;
        RECT 6.000 51.600 6.800 51.700 ;
        RECT 82.800 16.300 83.600 16.400 ;
        RECT 86.000 16.300 86.800 16.400 ;
        RECT 82.800 15.700 86.800 16.300 ;
        RECT 82.800 15.600 83.600 15.700 ;
        RECT 86.000 15.600 86.800 15.700 ;
    END
  END clk
  PIN in[1]
    PORT
      LAYER metal1 ;
        RECT 97.200 67.600 98.800 68.400 ;
        RECT 67.600 33.600 68.400 34.400 ;
        RECT 90.000 33.600 90.800 34.400 ;
        RECT 46.000 31.600 46.800 33.200 ;
        RECT 67.800 32.400 68.400 33.600 ;
        RECT 90.200 32.400 90.800 33.600 ;
        RECT 55.600 30.800 56.400 32.400 ;
        RECT 67.800 31.800 69.200 32.400 ;
        RECT 90.200 31.800 91.600 32.400 ;
        RECT 68.400 31.600 69.200 31.800 ;
        RECT 90.800 31.600 91.600 31.800 ;
        RECT 18.000 29.600 19.600 30.400 ;
        RECT 38.000 26.800 38.800 28.400 ;
        RECT 73.200 15.600 74.000 17.200 ;
        RECT 44.400 13.600 45.200 15.200 ;
      LAYER metal2 ;
        RECT 97.200 67.600 98.000 68.400 ;
        RECT 97.300 62.400 97.900 67.600 ;
        RECT 90.800 61.600 91.600 62.400 ;
        RECT 97.200 61.600 98.000 62.400 ;
        RECT 90.900 32.400 91.500 61.600 ;
        RECT 46.000 31.600 46.800 32.400 ;
        RECT 55.600 31.600 56.400 32.400 ;
        RECT 68.400 31.600 69.200 32.400 ;
        RECT 90.800 31.600 91.600 32.400 ;
        RECT 46.100 30.400 46.700 31.600 ;
        RECT 55.700 30.400 56.300 31.600 ;
        RECT 68.500 30.400 69.100 31.600 ;
        RECT 90.900 30.400 91.500 31.600 ;
        RECT 18.800 29.600 19.600 30.400 ;
        RECT 38.000 29.600 38.800 30.400 ;
        RECT 44.400 29.600 45.200 30.400 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 55.600 29.600 56.400 30.400 ;
        RECT 68.400 29.600 69.200 30.400 ;
        RECT 73.200 29.600 74.000 30.400 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 38.100 28.400 38.700 29.600 ;
        RECT 38.000 27.600 38.800 28.400 ;
        RECT 44.500 14.400 45.100 29.600 ;
        RECT 73.300 16.400 73.900 29.600 ;
        RECT 73.200 15.600 74.000 16.400 ;
        RECT 44.400 13.600 45.200 14.400 ;
        RECT 97.300 -2.300 97.900 29.600 ;
      LAYER metal3 ;
        RECT 90.800 62.300 91.600 62.400 ;
        RECT 97.200 62.300 98.000 62.400 ;
        RECT 90.800 61.700 98.000 62.300 ;
        RECT 90.800 61.600 91.600 61.700 ;
        RECT 97.200 61.600 98.000 61.700 ;
        RECT 18.800 30.300 19.600 30.400 ;
        RECT 38.000 30.300 38.800 30.400 ;
        RECT 44.400 30.300 45.200 30.400 ;
        RECT 46.000 30.300 46.800 30.400 ;
        RECT 55.600 30.300 56.400 30.400 ;
        RECT 68.400 30.300 69.200 30.400 ;
        RECT 73.200 30.300 74.000 30.400 ;
        RECT 90.800 30.300 91.600 30.400 ;
        RECT 97.200 30.300 98.000 30.400 ;
        RECT 18.800 29.700 98.000 30.300 ;
        RECT 18.800 29.600 19.600 29.700 ;
        RECT 38.000 29.600 38.800 29.700 ;
        RECT 44.400 29.600 45.200 29.700 ;
        RECT 46.000 29.600 46.800 29.700 ;
        RECT 55.600 29.600 56.400 29.700 ;
        RECT 68.400 29.600 69.200 29.700 ;
        RECT 73.200 29.600 74.000 29.700 ;
        RECT 90.800 29.600 91.600 29.700 ;
        RECT 97.200 29.600 98.000 29.700 ;
    END
  END in[1]
  PIN in[0]
    PORT
      LAYER metal1 ;
        RECT 100.000 67.600 100.800 68.400 ;
        RECT 106.000 68.300 107.600 68.400 ;
        RECT 110.000 68.300 110.800 68.400 ;
        RECT 106.000 68.200 110.800 68.300 ;
        RECT 100.200 67.200 100.800 67.600 ;
        RECT 104.200 67.700 110.800 68.200 ;
        RECT 104.200 67.600 107.600 67.700 ;
        RECT 110.000 67.600 110.800 67.700 ;
        RECT 104.200 67.200 104.800 67.600 ;
        RECT 100.200 66.400 101.000 67.200 ;
        RECT 102.800 66.600 104.800 67.200 ;
        RECT 102.800 66.400 104.400 66.600 ;
        RECT 58.000 33.600 58.800 34.400 ;
        RECT 58.000 32.400 58.600 33.600 ;
        RECT 57.200 31.800 58.600 32.400 ;
        RECT 57.200 31.600 58.000 31.800 ;
        RECT 49.200 26.800 50.000 28.400 ;
        RECT 42.800 24.800 43.600 26.400 ;
        RECT 64.400 14.400 65.200 14.800 ;
        RECT 64.400 13.800 66.000 14.400 ;
        RECT 65.200 13.600 66.000 13.800 ;
        RECT 70.000 13.600 70.800 15.200 ;
      LAYER metal2 ;
        RECT 110.000 67.600 110.800 68.400 ;
        RECT 100.200 67.000 101.000 67.200 ;
        RECT 103.600 67.000 104.400 67.200 ;
        RECT 100.200 66.400 104.400 67.000 ;
        RECT 49.200 31.600 50.000 32.400 ;
        RECT 57.200 32.300 58.000 32.400 ;
        RECT 57.200 31.700 59.500 32.300 ;
        RECT 57.200 31.600 58.000 31.700 ;
        RECT 49.300 28.400 49.900 31.600 ;
        RECT 49.200 27.600 50.000 28.400 ;
        RECT 49.300 26.400 49.900 27.600 ;
        RECT 42.800 25.600 43.600 26.400 ;
        RECT 49.200 25.600 50.000 26.400 ;
        RECT 58.900 14.400 59.500 31.700 ;
        RECT 110.100 14.400 110.700 67.600 ;
        RECT 58.800 13.600 59.600 14.400 ;
        RECT 65.200 13.600 66.000 14.400 ;
        RECT 70.000 13.600 70.800 14.400 ;
        RECT 110.000 13.600 110.800 14.400 ;
      LAYER metal3 ;
        RECT 110.000 68.300 110.800 68.400 ;
        RECT 110.000 67.700 113.900 68.300 ;
        RECT 110.000 67.600 110.800 67.700 ;
        RECT 49.200 32.300 50.000 32.400 ;
        RECT 57.200 32.300 58.000 32.400 ;
        RECT 49.200 31.700 58.000 32.300 ;
        RECT 49.200 31.600 50.000 31.700 ;
        RECT 57.200 31.600 58.000 31.700 ;
        RECT 42.800 26.300 43.600 26.400 ;
        RECT 49.200 26.300 50.000 26.400 ;
        RECT 42.800 25.700 50.000 26.300 ;
        RECT 42.800 25.600 43.600 25.700 ;
        RECT 49.200 25.600 50.000 25.700 ;
        RECT 58.800 14.300 59.600 14.400 ;
        RECT 65.200 14.300 66.000 14.400 ;
        RECT 70.000 14.300 70.800 14.400 ;
        RECT 110.000 14.300 110.800 14.400 ;
        RECT 58.800 13.700 110.800 14.300 ;
        RECT 58.800 13.600 59.600 13.700 ;
        RECT 65.200 13.600 66.000 13.700 ;
        RECT 70.000 13.600 70.800 13.700 ;
        RECT 110.000 13.600 110.800 13.700 ;
    END
  END in[0]
  PIN out
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER metal2 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 1.300 8.400 1.900 9.600 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -3.500 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END out
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 27.600 67.600 29.200 68.400 ;
        RECT 66.000 67.600 67.600 68.400 ;
        RECT 49.200 66.300 50.000 66.400 ;
        RECT 51.400 66.300 53.200 66.400 ;
        RECT 49.200 65.700 53.200 66.300 ;
        RECT 49.200 65.600 50.000 65.700 ;
        RECT 51.400 65.600 53.200 65.700 ;
        RECT 49.200 55.600 50.000 57.200 ;
        RECT 52.400 56.300 53.200 56.400 ;
        RECT 55.600 56.300 57.400 56.400 ;
        RECT 52.400 55.700 57.400 56.300 ;
        RECT 52.400 55.600 53.200 55.700 ;
        RECT 55.600 55.600 57.400 55.700 ;
        RECT 86.000 55.600 86.800 57.200 ;
        RECT 62.000 28.300 62.800 28.400 ;
        RECT 63.600 28.300 64.400 28.400 ;
        RECT 62.000 28.200 64.400 28.300 ;
        RECT 86.000 28.200 86.800 28.400 ;
        RECT 61.200 27.700 65.200 28.200 ;
        RECT 61.200 27.600 62.800 27.700 ;
        RECT 63.600 27.600 65.200 27.700 ;
        RECT 86.000 27.600 87.600 28.200 ;
        RECT 61.200 27.200 62.000 27.600 ;
        RECT 64.400 27.200 65.200 27.600 ;
        RECT 86.800 27.200 87.600 27.600 ;
      LAYER metal2 ;
        RECT 66.900 68.400 67.500 86.300 ;
        RECT 28.400 67.600 29.200 68.400 ;
        RECT 52.400 67.600 53.200 68.400 ;
        RECT 66.800 67.600 67.600 68.400 ;
        RECT 86.000 67.600 86.800 68.400 ;
        RECT 52.500 66.400 53.100 67.600 ;
        RECT 49.200 65.600 50.000 66.400 ;
        RECT 52.400 65.600 53.200 66.400 ;
        RECT 49.300 56.400 49.900 65.600 ;
        RECT 52.500 56.400 53.100 65.600 ;
        RECT 86.100 56.400 86.700 67.600 ;
        RECT 49.200 55.600 50.000 56.400 ;
        RECT 52.400 55.600 53.200 56.400 ;
        RECT 86.000 55.600 86.800 56.400 ;
        RECT 86.100 40.400 86.700 55.600 ;
        RECT 63.600 39.600 64.400 40.400 ;
        RECT 86.000 39.600 86.800 40.400 ;
        RECT 63.700 28.400 64.300 39.600 ;
        RECT 86.100 28.400 86.700 39.600 ;
        RECT 63.600 27.600 64.400 28.400 ;
        RECT 86.000 27.600 86.800 28.400 ;
      LAYER metal3 ;
        RECT 28.400 68.300 29.200 68.400 ;
        RECT 52.400 68.300 53.200 68.400 ;
        RECT 66.800 68.300 67.600 68.400 ;
        RECT 86.000 68.300 86.800 68.400 ;
        RECT 28.400 67.700 86.800 68.300 ;
        RECT 28.400 67.600 29.200 67.700 ;
        RECT 52.400 67.600 53.200 67.700 ;
        RECT 66.800 67.600 67.600 67.700 ;
        RECT 86.000 67.600 86.800 67.700 ;
        RECT 63.600 40.300 64.400 40.400 ;
        RECT 86.000 40.300 86.800 40.400 ;
        RECT 63.600 39.700 86.800 40.300 ;
        RECT 63.600 39.600 64.400 39.700 ;
        RECT 86.000 39.600 86.800 39.700 ;
    END
  END rst
  OBS
      LAYER metal1 ;
        RECT 1.200 71.400 2.000 79.800 ;
        RECT 5.600 76.400 6.400 79.800 ;
        RECT 4.400 75.800 6.400 76.400 ;
        RECT 10.000 75.800 10.800 79.800 ;
        RECT 14.200 75.800 15.400 79.800 ;
        RECT 4.400 75.000 5.200 75.800 ;
        RECT 10.000 75.200 10.600 75.800 ;
        RECT 7.800 74.600 11.400 75.200 ;
        RECT 14.000 75.000 14.800 75.800 ;
        RECT 7.800 74.400 8.600 74.600 ;
        RECT 10.600 74.400 11.400 74.600 ;
        RECT 4.400 73.000 5.200 73.200 ;
        RECT 9.000 73.000 9.800 73.200 ;
        RECT 4.400 72.400 9.800 73.000 ;
        RECT 10.400 73.000 12.600 73.600 ;
        RECT 10.400 71.800 11.000 73.000 ;
        RECT 11.800 72.800 12.600 73.000 ;
        RECT 6.200 71.400 11.000 71.800 ;
        RECT 1.200 71.200 11.000 71.400 ;
        RECT 18.800 71.200 19.600 79.800 ;
        RECT 20.600 79.200 24.200 79.800 ;
        RECT 20.600 79.000 21.200 79.200 ;
        RECT 20.400 73.000 21.200 79.000 ;
        RECT 23.600 79.000 24.200 79.200 ;
        RECT 25.200 79.200 29.200 79.800 ;
        RECT 22.000 73.000 22.800 78.600 ;
        RECT 23.600 73.400 24.400 79.000 ;
        RECT 25.200 74.000 26.000 79.200 ;
        RECT 26.800 73.800 27.600 78.600 ;
        RECT 28.400 73.800 29.200 79.200 ;
        RECT 26.800 73.400 27.400 73.800 ;
        RECT 23.600 73.000 27.400 73.400 ;
        RECT 22.200 72.400 22.800 73.000 ;
        RECT 23.800 72.800 27.400 73.000 ;
        RECT 28.600 73.200 29.200 73.800 ;
        RECT 31.600 73.800 32.400 79.800 ;
        RECT 31.600 73.200 32.200 73.800 ;
        RECT 28.600 72.600 32.200 73.200 ;
        RECT 22.000 72.200 22.800 72.400 ;
        RECT 22.000 71.600 25.400 72.200 ;
        RECT 1.200 71.000 7.000 71.200 ;
        RECT 1.200 70.800 6.800 71.000 ;
        RECT 15.400 70.600 19.600 71.200 ;
        RECT 15.400 70.400 16.200 70.600 ;
        RECT 7.600 70.200 8.400 70.400 ;
        RECT 3.400 69.600 8.400 70.200 ;
        RECT 17.000 69.800 17.800 70.000 ;
        RECT 3.400 69.400 4.200 69.600 ;
        RECT 14.000 69.200 17.800 69.800 ;
        RECT 14.000 69.000 14.800 69.200 ;
        RECT 18.800 67.200 19.600 70.600 ;
        RECT 1.200 62.200 2.000 67.000 ;
        RECT 15.800 66.600 19.600 67.200 ;
        RECT 15.800 66.400 16.600 66.600 ;
        RECT 7.800 65.400 8.600 65.600 ;
        RECT 4.400 64.200 5.200 65.000 ;
        RECT 7.800 64.800 10.600 65.400 ;
        RECT 10.000 64.200 10.600 64.800 ;
        RECT 14.000 64.200 14.800 65.000 ;
        RECT 4.400 63.600 6.400 64.200 ;
        RECT 5.600 62.200 6.400 63.600 ;
        RECT 10.000 62.200 10.800 64.200 ;
        RECT 14.000 63.600 15.400 64.200 ;
        RECT 14.200 62.200 15.400 63.600 ;
        RECT 18.800 62.200 19.600 66.600 ;
        RECT 24.800 65.000 25.400 71.600 ;
        RECT 26.000 70.300 27.600 70.400 ;
        RECT 39.600 70.300 40.400 79.800 ;
        RECT 43.000 79.200 46.600 79.800 ;
        RECT 43.000 79.000 43.600 79.200 ;
        RECT 42.800 73.000 43.600 79.000 ;
        RECT 46.000 79.000 46.600 79.200 ;
        RECT 47.600 79.200 51.600 79.800 ;
        RECT 44.400 73.000 45.200 78.600 ;
        RECT 46.000 73.400 46.800 79.000 ;
        RECT 47.600 74.000 48.400 79.200 ;
        RECT 49.200 73.800 50.000 78.600 ;
        RECT 50.800 73.800 51.600 79.200 ;
        RECT 49.200 73.400 49.800 73.800 ;
        RECT 46.000 73.000 49.800 73.400 ;
        RECT 44.600 72.400 45.200 73.000 ;
        RECT 46.200 72.800 49.800 73.000 ;
        RECT 51.000 73.200 51.600 73.800 ;
        RECT 54.000 73.800 54.800 79.800 ;
        RECT 54.000 73.200 54.600 73.800 ;
        RECT 51.000 72.600 54.600 73.200 ;
        RECT 44.400 72.200 45.200 72.400 ;
        RECT 44.400 71.600 47.800 72.200 ;
        RECT 44.400 70.300 45.200 70.400 ;
        RECT 26.000 69.700 45.200 70.300 ;
        RECT 26.000 69.600 27.600 69.700 ;
        RECT 29.000 65.600 30.800 66.400 ;
        RECT 24.800 64.400 28.800 65.000 ;
        RECT 20.400 64.300 21.200 64.400 ;
        RECT 24.800 64.300 26.000 64.400 ;
        RECT 20.400 63.700 26.000 64.300 ;
        RECT 20.400 63.600 21.200 63.700 ;
        RECT 25.200 62.200 26.000 63.700 ;
        RECT 28.200 64.200 28.800 64.400 ;
        RECT 28.200 63.600 29.200 64.200 ;
        RECT 28.400 62.200 29.200 63.600 ;
        RECT 39.600 62.200 40.400 69.700 ;
        RECT 44.400 69.600 45.200 69.700 ;
        RECT 41.200 66.300 42.000 66.400 ;
        RECT 42.800 66.300 43.600 66.400 ;
        RECT 41.200 65.700 43.600 66.300 ;
        RECT 41.200 64.800 42.000 65.700 ;
        RECT 42.800 65.600 43.600 65.700 ;
        RECT 47.200 65.000 47.800 71.600 ;
        RECT 48.400 69.600 50.000 70.400 ;
        RECT 50.000 68.300 51.600 68.400 ;
        RECT 57.200 68.300 58.000 79.800 ;
        RECT 59.000 79.200 62.600 79.800 ;
        RECT 59.000 79.000 59.600 79.200 ;
        RECT 58.800 73.000 59.600 79.000 ;
        RECT 62.000 79.000 62.600 79.200 ;
        RECT 63.600 79.200 67.600 79.800 ;
        RECT 60.400 73.000 61.200 78.600 ;
        RECT 62.000 73.400 62.800 79.000 ;
        RECT 63.600 74.000 64.400 79.200 ;
        RECT 65.200 73.800 66.000 78.600 ;
        RECT 66.800 73.800 67.600 79.200 ;
        RECT 65.200 73.400 65.800 73.800 ;
        RECT 62.000 73.000 65.800 73.400 ;
        RECT 60.600 72.400 61.200 73.000 ;
        RECT 62.200 72.800 65.800 73.000 ;
        RECT 67.000 73.200 67.600 73.800 ;
        RECT 70.000 73.800 70.800 79.800 ;
        RECT 70.000 73.200 70.600 73.800 ;
        RECT 67.000 72.600 70.600 73.200 ;
        RECT 60.400 72.200 61.200 72.400 ;
        RECT 60.400 71.600 63.800 72.200 ;
        RECT 50.000 67.700 58.000 68.300 ;
        RECT 50.000 67.600 51.600 67.700 ;
        RECT 47.200 64.400 51.200 65.000 ;
        RECT 55.600 64.800 56.400 66.400 ;
        RECT 47.200 64.200 48.400 64.400 ;
        RECT 47.600 62.200 48.400 64.200 ;
        RECT 50.600 63.600 51.600 64.400 ;
        RECT 50.800 62.200 51.600 63.600 ;
        RECT 57.200 64.300 58.000 67.700 ;
        RECT 63.200 65.000 63.800 71.600 ;
        RECT 78.000 71.400 78.800 79.800 ;
        RECT 82.400 76.400 83.200 79.800 ;
        RECT 81.200 75.800 83.200 76.400 ;
        RECT 86.800 75.800 87.600 79.800 ;
        RECT 91.000 75.800 92.200 79.800 ;
        RECT 81.200 75.000 82.000 75.800 ;
        RECT 86.800 75.200 87.400 75.800 ;
        RECT 84.600 74.600 88.200 75.200 ;
        RECT 90.800 75.000 91.600 75.800 ;
        RECT 84.600 74.400 85.400 74.600 ;
        RECT 87.400 74.400 88.200 74.600 ;
        RECT 81.200 73.000 82.000 73.200 ;
        RECT 85.800 73.000 86.600 73.200 ;
        RECT 81.200 72.400 86.600 73.000 ;
        RECT 87.200 73.000 89.400 73.600 ;
        RECT 87.200 71.800 87.800 73.000 ;
        RECT 88.600 72.800 89.400 73.000 ;
        RECT 83.000 71.400 87.800 71.800 ;
        RECT 78.000 71.200 87.800 71.400 ;
        RECT 95.600 71.200 96.400 79.800 ;
        RECT 97.200 72.400 98.000 79.800 ;
        RECT 98.800 72.400 99.600 72.600 ;
        RECT 101.600 72.400 103.200 79.800 ;
        RECT 97.200 71.800 99.600 72.400 ;
        RECT 101.200 71.800 103.200 72.400 ;
        RECT 105.400 72.400 106.200 72.600 ;
        RECT 106.800 72.400 107.600 79.800 ;
        RECT 105.400 71.800 107.600 72.400 ;
        RECT 78.000 71.000 83.800 71.200 ;
        RECT 78.000 70.800 83.600 71.000 ;
        RECT 92.200 70.600 96.400 71.200 ;
        RECT 92.200 70.400 93.000 70.600 ;
        RECT 64.400 69.600 66.000 70.400 ;
        RECT 84.400 70.200 85.200 70.400 ;
        RECT 80.200 69.600 85.200 70.200 ;
        RECT 93.800 69.800 94.600 70.000 ;
        RECT 80.200 69.400 81.000 69.600 ;
        RECT 90.800 69.200 94.600 69.800 ;
        RECT 90.800 69.000 91.600 69.200 ;
        RECT 95.600 67.200 96.400 70.600 ;
        RECT 101.200 70.400 101.800 71.800 ;
        RECT 105.400 71.200 106.000 71.800 ;
        RECT 102.600 70.600 106.000 71.200 ;
        RECT 102.600 70.400 103.400 70.600 ;
        RECT 100.400 69.800 101.800 70.400 ;
        RECT 104.800 69.800 105.600 70.000 ;
        RECT 100.400 69.600 102.200 69.800 ;
        RECT 101.200 69.200 102.200 69.600 ;
        RECT 66.800 65.600 69.200 66.400 ;
        RECT 63.200 64.400 67.200 65.000 ;
        RECT 58.800 64.300 59.600 64.400 ;
        RECT 57.200 63.700 59.600 64.300 ;
        RECT 63.200 64.200 64.400 64.400 ;
        RECT 57.200 62.200 58.000 63.700 ;
        RECT 58.800 63.600 59.600 63.700 ;
        RECT 63.600 62.200 64.400 64.200 ;
        RECT 66.600 64.200 67.200 64.400 ;
        RECT 66.600 63.600 67.600 64.200 ;
        RECT 66.800 62.200 67.600 63.600 ;
        RECT 78.000 62.200 78.800 67.000 ;
        RECT 92.600 66.600 96.400 67.200 ;
        RECT 98.800 66.800 99.600 67.000 ;
        RECT 92.600 66.400 93.400 66.600 ;
        RECT 84.600 65.400 85.400 65.600 ;
        RECT 81.200 64.200 82.000 65.000 ;
        RECT 84.600 64.800 87.400 65.400 ;
        RECT 86.800 64.200 87.400 64.800 ;
        RECT 90.800 64.200 91.600 65.000 ;
        RECT 81.200 63.600 83.200 64.200 ;
        RECT 82.400 62.200 83.200 63.600 ;
        RECT 86.800 62.200 87.600 64.200 ;
        RECT 90.800 63.600 92.200 64.200 ;
        RECT 91.000 62.200 92.200 63.600 ;
        RECT 95.600 62.200 96.400 66.600 ;
        RECT 97.200 66.200 99.600 66.800 ;
        RECT 97.200 62.200 98.000 66.200 ;
        RECT 101.600 65.800 102.200 69.200 ;
        RECT 103.000 69.200 105.600 69.800 ;
        RECT 103.000 68.600 103.600 69.200 ;
        RECT 102.800 67.800 103.600 68.600 ;
        RECT 105.400 66.800 106.200 67.000 ;
        RECT 105.400 66.200 107.600 66.800 ;
        RECT 101.600 64.400 103.200 65.800 ;
        RECT 100.400 63.600 103.200 64.400 ;
        RECT 101.600 62.200 103.200 63.600 ;
        RECT 106.800 62.200 107.600 66.200 ;
        RECT 1.200 55.000 2.000 59.800 ;
        RECT 5.600 58.400 6.400 59.800 ;
        RECT 4.400 57.800 6.400 58.400 ;
        RECT 10.000 57.800 10.800 59.800 ;
        RECT 14.200 58.400 15.400 59.800 ;
        RECT 14.000 57.800 15.400 58.400 ;
        RECT 4.400 57.000 5.200 57.800 ;
        RECT 10.000 57.200 10.600 57.800 ;
        RECT 7.800 56.600 10.600 57.200 ;
        RECT 14.000 57.000 14.800 57.800 ;
        RECT 7.800 56.400 8.600 56.600 ;
        RECT 15.800 55.400 16.600 55.600 ;
        RECT 18.800 55.400 19.600 59.800 ;
        RECT 20.400 56.000 21.200 59.800 ;
        RECT 23.600 56.000 24.400 59.800 ;
        RECT 20.400 55.800 24.400 56.000 ;
        RECT 25.200 55.800 26.000 59.800 ;
        RECT 33.800 56.400 34.600 59.800 ;
        RECT 38.600 58.400 39.400 59.800 ;
        RECT 38.000 57.600 39.400 58.400 ;
        RECT 38.600 56.400 39.400 57.600 ;
        RECT 33.800 55.800 35.600 56.400 ;
        RECT 38.600 55.800 40.400 56.400 ;
        RECT 42.800 56.000 43.600 59.800 ;
        RECT 46.000 56.000 46.800 59.800 ;
        RECT 42.800 55.800 46.800 56.000 ;
        RECT 47.600 55.800 48.400 59.800 ;
        RECT 50.800 57.800 51.600 59.800 ;
        RECT 57.200 58.400 58.000 59.800 ;
        RECT 57.200 57.800 58.200 58.400 ;
        RECT 20.600 55.400 24.200 55.800 ;
        RECT 15.800 54.800 19.600 55.400 ;
        RECT 18.800 54.300 19.600 54.800 ;
        RECT 21.200 54.400 22.000 54.800 ;
        RECT 25.200 54.400 25.800 55.800 ;
        RECT 20.400 54.300 22.000 54.400 ;
        RECT 18.800 53.800 22.000 54.300 ;
        RECT 18.800 53.700 21.200 53.800 ;
        RECT 14.000 52.800 14.800 53.000 ;
        RECT 3.400 52.400 4.200 52.600 ;
        RECT 3.400 51.800 8.400 52.400 ;
        RECT 14.000 52.200 17.800 52.800 ;
        RECT 17.000 52.000 17.800 52.200 ;
        RECT 7.600 51.600 8.400 51.800 ;
        RECT 15.400 51.400 16.200 51.600 ;
        RECT 18.800 51.400 19.600 53.700 ;
        RECT 20.400 53.600 21.200 53.700 ;
        RECT 23.400 53.600 26.000 54.400 ;
        RECT 22.000 51.600 22.800 53.200 ;
        RECT 23.400 52.400 24.000 53.600 ;
        RECT 23.400 51.600 24.400 52.400 ;
        RECT 1.200 51.000 6.800 51.200 ;
        RECT 1.200 50.800 7.000 51.000 ;
        RECT 15.400 50.800 19.600 51.400 ;
        RECT 1.200 50.600 11.000 50.800 ;
        RECT 1.200 42.200 2.000 50.600 ;
        RECT 6.200 50.200 11.000 50.600 ;
        RECT 4.400 49.000 9.800 49.600 ;
        RECT 4.400 48.800 5.200 49.000 ;
        RECT 9.000 48.800 9.800 49.000 ;
        RECT 10.400 49.000 11.000 50.200 ;
        RECT 11.800 49.000 12.600 49.200 ;
        RECT 10.400 48.400 12.600 49.000 ;
        RECT 7.800 47.400 8.600 47.600 ;
        RECT 10.600 47.400 11.400 47.600 ;
        RECT 4.400 46.200 5.200 47.000 ;
        RECT 7.800 46.800 11.400 47.400 ;
        RECT 10.000 46.200 10.600 46.800 ;
        RECT 14.000 46.200 14.800 47.000 ;
        RECT 4.400 45.600 6.400 46.200 ;
        RECT 5.600 42.200 6.400 45.600 ;
        RECT 10.000 42.200 10.800 46.200 ;
        RECT 14.200 42.200 15.400 46.200 ;
        RECT 18.800 42.200 19.600 50.800 ;
        RECT 23.400 50.200 24.000 51.600 ;
        RECT 25.200 50.200 26.000 50.400 ;
        RECT 23.000 49.600 24.000 50.200 ;
        RECT 24.600 49.600 26.000 50.200 ;
        RECT 23.000 42.200 23.800 49.600 ;
        RECT 24.600 48.400 25.200 49.600 ;
        RECT 33.200 48.800 34.000 50.400 ;
        RECT 34.800 50.300 35.600 55.800 ;
        RECT 36.400 53.600 37.200 55.200 ;
        RECT 38.000 50.300 38.800 50.400 ;
        RECT 34.800 49.700 38.800 50.300 ;
        RECT 24.400 47.600 25.200 48.400 ;
        RECT 34.800 42.200 35.600 49.700 ;
        RECT 38.000 48.800 38.800 49.700 ;
        RECT 39.600 42.200 40.400 55.800 ;
        RECT 43.000 55.400 46.600 55.800 ;
        RECT 41.200 53.600 42.000 55.200 ;
        RECT 43.600 54.400 44.400 54.800 ;
        RECT 47.600 54.400 48.200 55.800 ;
        RECT 51.000 54.400 51.600 57.800 ;
        RECT 57.600 57.600 58.200 57.800 ;
        RECT 60.400 57.800 61.200 59.800 ;
        RECT 60.400 57.600 61.600 57.800 ;
        RECT 57.600 57.000 61.600 57.600 ;
        RECT 61.000 54.400 61.600 57.000 ;
        RECT 66.800 56.000 67.600 59.800 ;
        RECT 70.000 56.000 70.800 59.800 ;
        RECT 66.800 55.800 70.800 56.000 ;
        RECT 71.600 55.800 72.400 59.800 ;
        RECT 73.400 56.400 74.200 57.200 ;
        RECT 67.000 55.400 70.600 55.800 ;
        RECT 67.600 54.400 68.400 54.800 ;
        RECT 71.600 54.400 72.200 55.800 ;
        RECT 73.200 55.600 74.000 56.400 ;
        RECT 74.800 55.800 75.600 59.800 ;
        RECT 42.800 53.800 44.400 54.400 ;
        RECT 42.800 53.600 43.600 53.800 ;
        RECT 45.800 53.600 48.400 54.400 ;
        RECT 50.800 53.600 51.600 54.400 ;
        RECT 57.200 53.600 58.800 54.400 ;
        RECT 60.400 53.600 61.600 54.400 ;
        RECT 66.800 53.800 68.400 54.400 ;
        RECT 66.800 53.600 67.600 53.800 ;
        RECT 69.800 53.600 72.400 54.400 ;
        RECT 44.400 51.600 45.200 53.200 ;
        RECT 45.800 50.200 46.400 53.600 ;
        RECT 51.000 52.300 51.600 53.600 ;
        RECT 47.700 51.700 51.600 52.300 ;
        RECT 47.700 50.400 48.300 51.700 ;
        RECT 47.600 50.200 48.400 50.400 ;
        RECT 51.000 50.200 51.600 51.700 ;
        RECT 52.400 52.300 53.200 52.400 ;
        RECT 58.800 52.300 60.400 52.400 ;
        RECT 52.400 51.700 60.400 52.300 ;
        RECT 52.400 50.800 53.200 51.700 ;
        RECT 58.800 51.600 60.400 51.700 ;
        RECT 61.000 50.400 61.600 53.600 ;
        RECT 68.400 51.600 69.200 53.200 ;
        RECT 69.800 52.400 70.400 53.600 ;
        RECT 75.000 52.400 75.600 55.800 ;
        RECT 76.400 52.800 77.200 54.400 ;
        RECT 69.800 51.600 70.800 52.400 ;
        RECT 73.200 52.200 74.000 52.400 ;
        RECT 74.800 52.200 75.600 52.400 ;
        RECT 78.000 52.300 78.800 52.400 ;
        RECT 87.600 52.300 88.400 59.800 ;
        RECT 92.400 55.800 93.200 59.800 ;
        RECT 93.800 56.400 94.600 57.200 ;
        RECT 89.200 54.300 90.000 54.400 ;
        RECT 90.800 54.300 91.600 54.400 ;
        RECT 89.200 53.700 91.600 54.300 ;
        RECT 89.200 53.600 90.000 53.700 ;
        RECT 90.800 52.800 91.600 53.700 ;
        RECT 89.200 52.300 90.000 52.400 ;
        RECT 78.000 52.200 90.000 52.300 ;
        RECT 92.400 52.200 93.000 55.800 ;
        RECT 94.000 55.600 94.800 56.400 ;
        RECT 98.600 55.800 100.200 59.800 ;
        RECT 97.200 52.800 98.000 54.400 ;
        RECT 99.000 52.400 99.600 55.800 ;
        RECT 100.400 53.600 101.200 54.400 ;
        RECT 107.200 54.200 108.000 59.800 ;
        RECT 107.200 53.800 109.000 54.200 ;
        RECT 107.400 53.600 109.000 53.800 ;
        RECT 100.400 53.200 101.000 53.600 ;
        RECT 100.200 52.400 101.000 53.200 ;
        RECT 94.000 52.200 94.800 52.400 ;
        RECT 73.200 51.600 75.600 52.200 ;
        RECT 77.200 51.700 90.800 52.200 ;
        RECT 77.200 51.600 78.800 51.700 ;
        RECT 45.400 49.600 46.400 50.200 ;
        RECT 47.000 49.600 48.400 50.200 ;
        RECT 45.400 42.200 46.200 49.600 ;
        RECT 47.000 48.400 47.600 49.600 ;
        RECT 50.800 49.400 52.600 50.200 ;
        RECT 61.000 49.800 64.400 50.400 ;
        RECT 69.800 50.200 70.400 51.600 ;
        RECT 71.600 50.200 72.400 50.400 ;
        RECT 73.400 50.200 74.000 51.600 ;
        RECT 77.200 51.200 78.000 51.600 ;
        RECT 63.600 49.600 64.400 49.800 ;
        RECT 69.400 49.600 70.400 50.200 ;
        RECT 71.000 49.600 72.400 50.200 ;
        RECT 46.800 47.600 47.600 48.400 ;
        RECT 51.800 42.200 52.600 49.400 ;
        RECT 54.200 48.800 57.800 49.400 ;
        RECT 54.200 48.200 54.800 48.800 ;
        RECT 54.000 42.200 54.800 48.200 ;
        RECT 57.200 48.200 57.800 48.800 ;
        RECT 59.000 49.000 62.600 49.200 ;
        RECT 63.600 49.000 64.200 49.600 ;
        RECT 59.000 48.600 62.800 49.000 ;
        RECT 59.000 48.200 59.600 48.600 ;
        RECT 57.200 42.800 58.000 48.200 ;
        RECT 58.800 43.400 59.600 48.200 ;
        RECT 60.400 42.800 61.200 48.000 ;
        RECT 62.000 43.000 62.800 48.600 ;
        RECT 63.600 43.400 64.400 49.000 ;
        RECT 57.200 42.200 61.200 42.800 ;
        RECT 62.200 42.800 62.800 43.000 ;
        RECT 65.200 43.000 66.000 49.000 ;
        RECT 65.200 42.800 65.800 43.000 ;
        RECT 62.200 42.200 65.800 42.800 ;
        RECT 69.400 42.200 70.200 49.600 ;
        RECT 71.000 48.400 71.600 49.600 ;
        RECT 70.800 47.600 71.600 48.400 ;
        RECT 73.200 42.200 74.000 50.200 ;
        RECT 74.800 49.600 78.800 50.200 ;
        RECT 74.800 42.200 75.600 49.600 ;
        RECT 78.000 42.200 78.800 49.600 ;
        RECT 87.600 42.200 88.400 51.700 ;
        RECT 89.200 51.600 90.800 51.700 ;
        RECT 92.400 51.600 94.800 52.200 ;
        RECT 95.600 52.200 96.400 52.400 ;
        RECT 95.600 51.600 97.200 52.200 ;
        RECT 98.800 51.600 99.600 52.400 ;
        RECT 90.000 51.200 90.800 51.600 ;
        RECT 94.000 50.200 94.600 51.600 ;
        RECT 96.400 51.200 97.200 51.600 ;
        RECT 99.000 51.400 99.600 51.600 ;
        RECT 99.000 50.800 101.000 51.400 ;
        RECT 102.000 50.800 102.800 52.400 ;
        RECT 105.200 51.600 106.800 52.400 ;
        RECT 100.400 50.200 101.000 50.800 ;
        RECT 89.200 49.600 93.200 50.200 ;
        RECT 89.200 42.200 90.000 49.600 ;
        RECT 92.400 42.200 93.200 49.600 ;
        RECT 94.000 42.200 94.800 50.200 ;
        RECT 95.600 49.600 99.600 50.200 ;
        RECT 95.600 42.200 96.400 49.600 ;
        RECT 98.800 42.800 99.600 49.600 ;
        RECT 100.400 43.400 101.200 50.200 ;
        RECT 102.000 42.800 102.800 50.200 ;
        RECT 103.600 49.600 104.400 51.200 ;
        RECT 108.400 50.400 109.000 53.600 ;
        RECT 108.400 49.600 109.200 50.400 ;
        RECT 106.800 47.600 107.600 49.200 ;
        RECT 108.400 47.000 109.000 49.600 ;
        RECT 105.400 46.400 109.000 47.000 ;
        RECT 98.800 42.200 102.800 42.800 ;
        RECT 105.200 42.200 106.000 46.400 ;
        RECT 108.400 46.200 109.000 46.400 ;
        RECT 108.400 42.200 109.200 46.200 ;
        RECT 1.200 35.800 2.000 39.800 ;
        RECT 1.400 35.600 2.000 35.800 ;
        RECT 4.400 35.800 5.200 39.800 ;
        RECT 4.400 35.600 5.000 35.800 ;
        RECT 1.400 35.000 5.000 35.600 ;
        RECT 1.400 32.400 2.000 35.000 ;
        RECT 2.800 32.800 3.600 34.400 ;
        RECT 1.200 31.600 2.000 32.400 ;
        RECT 1.400 28.400 2.000 31.600 ;
        RECT 6.000 30.800 6.800 32.400 ;
        RECT 7.600 31.600 8.400 33.200 ;
        RECT 3.600 29.600 5.200 30.400 ;
        RECT 7.600 30.300 8.400 30.400 ;
        RECT 9.200 30.300 10.000 39.800 ;
        RECT 7.600 29.700 10.000 30.300 ;
        RECT 7.600 29.600 8.400 29.700 ;
        RECT 1.400 28.200 3.000 28.400 ;
        RECT 1.400 27.800 3.200 28.200 ;
        RECT 2.400 22.200 3.200 27.800 ;
        RECT 9.200 26.200 10.000 29.700 ;
        RECT 12.400 32.300 13.200 39.800 ;
        RECT 15.600 35.800 16.400 39.800 ;
        RECT 15.800 35.600 16.400 35.800 ;
        RECT 18.800 35.800 19.600 39.800 ;
        RECT 18.800 35.600 19.400 35.800 ;
        RECT 15.800 35.000 19.400 35.600 ;
        RECT 14.000 34.300 14.800 34.400 ;
        RECT 15.800 34.300 16.400 35.000 ;
        RECT 14.000 33.700 16.400 34.300 ;
        RECT 14.000 33.600 14.800 33.700 ;
        RECT 15.800 32.400 16.400 33.700 ;
        RECT 17.200 32.800 18.000 34.400 ;
        RECT 14.000 32.300 14.800 32.400 ;
        RECT 12.400 31.700 14.800 32.300 ;
        RECT 10.800 28.300 11.600 28.400 ;
        RECT 12.400 28.300 13.200 31.700 ;
        RECT 14.000 31.600 14.800 31.700 ;
        RECT 15.600 31.600 16.400 32.400 ;
        RECT 10.800 27.700 13.200 28.300 ;
        RECT 15.800 28.400 16.400 31.600 ;
        RECT 20.400 30.800 21.200 32.400 ;
        RECT 15.800 28.200 17.400 28.400 ;
        RECT 15.800 27.800 17.600 28.200 ;
        RECT 10.800 26.800 11.600 27.700 ;
        RECT 8.200 25.600 10.000 26.200 ;
        RECT 8.200 22.200 9.000 25.600 ;
        RECT 12.400 22.200 13.200 27.700 ;
        RECT 14.000 24.800 14.800 26.400 ;
        RECT 16.800 22.200 17.600 27.800 ;
        RECT 22.000 22.200 22.800 39.800 ;
        RECT 25.200 32.400 26.000 39.800 ;
        RECT 28.400 32.400 29.200 39.800 ;
        RECT 25.200 31.800 29.200 32.400 ;
        RECT 30.000 31.800 30.800 39.800 ;
        RECT 26.000 30.400 26.800 30.800 ;
        RECT 30.000 30.400 30.600 31.800 ;
        RECT 25.200 29.800 26.800 30.400 ;
        RECT 28.400 29.800 30.800 30.400 ;
        RECT 25.200 29.600 26.000 29.800 ;
        RECT 26.800 27.600 27.600 29.200 ;
        RECT 23.600 24.800 24.400 26.400 ;
        RECT 28.400 26.200 29.000 29.800 ;
        RECT 30.000 29.600 30.800 29.800 ;
        RECT 28.400 22.200 29.200 26.200 ;
        RECT 30.000 25.600 30.800 26.400 ;
        RECT 39.600 26.200 40.400 39.800 ;
        RECT 41.200 32.300 42.000 34.400 ;
        RECT 44.400 32.300 45.200 39.800 ;
        RECT 41.200 31.700 45.200 32.300 ;
        RECT 41.200 31.600 42.000 31.700 ;
        RECT 39.600 25.600 41.400 26.200 ;
        RECT 29.800 24.800 30.600 25.600 ;
        RECT 40.600 24.400 41.400 25.600 ;
        RECT 40.600 23.600 42.000 24.400 ;
        RECT 40.600 22.200 41.400 23.600 ;
        RECT 44.400 22.200 45.200 31.700 ;
        RECT 46.000 28.300 46.800 28.400 ;
        RECT 47.600 28.300 48.400 39.800 ;
        RECT 50.800 35.800 51.600 39.800 ;
        RECT 51.000 35.600 51.600 35.800 ;
        RECT 54.000 35.800 54.800 39.800 ;
        RECT 54.000 35.600 54.600 35.800 ;
        RECT 51.000 35.000 54.600 35.600 ;
        RECT 51.000 32.400 51.600 35.000 ;
        RECT 52.400 32.800 53.200 34.400 ;
        RECT 59.400 32.400 60.200 39.800 ;
        RECT 50.800 31.600 51.600 32.400 ;
        RECT 46.000 27.700 48.400 28.300 ;
        RECT 51.000 28.400 51.600 31.600 ;
        RECT 59.200 31.800 60.200 32.400 ;
        RECT 66.200 32.400 67.000 39.800 ;
        RECT 71.600 35.800 72.400 39.800 ;
        RECT 71.800 35.600 72.400 35.800 ;
        RECT 74.800 38.300 75.600 39.800 ;
        RECT 81.200 38.300 82.000 38.400 ;
        RECT 74.800 37.700 82.000 38.300 ;
        RECT 74.800 35.800 75.600 37.700 ;
        RECT 81.200 37.600 82.000 37.700 ;
        RECT 76.400 36.300 77.200 36.400 ;
        RECT 82.800 36.300 83.600 39.800 ;
        RECT 74.800 35.600 75.400 35.800 ;
        RECT 76.400 35.700 83.600 36.300 ;
        RECT 76.400 35.600 77.200 35.700 ;
        RECT 71.800 35.000 75.400 35.600 ;
        RECT 73.200 32.800 74.000 34.400 ;
        RECT 74.800 32.400 75.400 35.000 ;
        RECT 66.200 31.800 67.200 32.400 ;
        RECT 53.200 29.600 54.800 30.400 ;
        RECT 59.200 28.400 59.800 31.800 ;
        RECT 60.400 30.300 61.200 30.400 ;
        RECT 65.200 30.300 66.000 30.400 ;
        RECT 60.400 29.700 66.000 30.300 ;
        RECT 60.400 28.800 61.200 29.700 ;
        RECT 65.200 28.800 66.000 29.700 ;
        RECT 51.000 28.200 52.600 28.400 ;
        RECT 51.000 27.800 52.800 28.200 ;
        RECT 46.000 27.600 46.800 27.700 ;
        RECT 47.600 26.200 48.400 27.700 ;
        RECT 46.600 25.600 48.400 26.200 ;
        RECT 46.600 22.200 47.400 25.600 ;
        RECT 52.000 22.200 52.800 27.800 ;
        RECT 57.200 27.600 59.800 28.400 ;
        RECT 66.600 28.400 67.200 31.800 ;
        RECT 70.000 30.800 70.800 32.400 ;
        RECT 74.800 31.600 75.600 32.400 ;
        RECT 71.600 29.600 73.200 30.400 ;
        RECT 74.800 28.400 75.400 31.600 ;
        RECT 66.600 27.600 69.200 28.400 ;
        RECT 73.800 28.200 75.400 28.400 ;
        RECT 73.600 27.800 75.400 28.200 ;
        RECT 57.400 26.200 58.000 27.600 ;
        RECT 59.000 26.200 62.600 26.600 ;
        RECT 63.800 26.200 67.400 26.600 ;
        RECT 68.400 26.200 69.000 27.600 ;
        RECT 57.200 22.200 58.000 26.200 ;
        RECT 58.800 26.000 62.800 26.200 ;
        RECT 58.800 22.200 59.600 26.000 ;
        RECT 62.000 22.200 62.800 26.000 ;
        RECT 63.600 26.000 67.600 26.200 ;
        RECT 63.600 22.200 64.400 26.000 ;
        RECT 66.800 22.200 67.600 26.000 ;
        RECT 68.400 22.200 69.200 26.200 ;
        RECT 73.600 22.200 74.400 27.800 ;
        RECT 82.800 22.200 83.600 35.700 ;
        RECT 88.600 32.400 89.400 39.800 ;
        RECT 94.000 35.800 94.800 39.800 ;
        RECT 94.200 35.600 94.800 35.800 ;
        RECT 97.200 35.800 98.000 39.800 ;
        RECT 97.200 35.600 97.800 35.800 ;
        RECT 94.200 35.000 97.800 35.600 ;
        RECT 95.600 32.800 96.400 34.400 ;
        RECT 97.200 32.400 97.800 35.000 ;
        RECT 98.800 32.400 99.600 39.800 ;
        RECT 105.800 38.400 106.600 39.800 ;
        RECT 105.800 37.600 107.600 38.400 ;
        RECT 104.400 33.600 105.200 34.400 ;
        RECT 104.400 32.400 105.000 33.600 ;
        RECT 105.800 32.400 106.600 37.600 ;
        RECT 88.600 31.800 89.600 32.400 ;
        RECT 87.600 28.800 88.400 30.400 ;
        RECT 89.000 28.400 89.600 31.800 ;
        RECT 92.400 30.800 93.200 32.400 ;
        RECT 97.200 31.600 98.000 32.400 ;
        RECT 98.800 31.800 101.000 32.400 ;
        RECT 94.000 29.600 95.600 30.400 ;
        RECT 97.200 28.400 97.800 31.600 ;
        RECT 100.400 31.200 101.000 31.800 ;
        RECT 103.600 31.800 105.000 32.400 ;
        RECT 105.600 31.800 106.600 32.400 ;
        RECT 103.600 31.600 104.400 31.800 ;
        RECT 100.400 30.400 101.600 31.200 ;
        RECT 98.800 28.800 99.600 30.400 ;
        RECT 89.000 27.600 91.600 28.400 ;
        RECT 96.200 28.200 97.800 28.400 ;
        RECT 96.000 27.800 97.800 28.200 ;
        RECT 84.400 24.800 85.200 26.400 ;
        RECT 86.200 26.200 89.800 26.600 ;
        RECT 90.800 26.200 91.400 27.600 ;
        RECT 86.000 26.000 90.000 26.200 ;
        RECT 86.000 22.200 86.800 26.000 ;
        RECT 89.200 22.200 90.000 26.000 ;
        RECT 90.800 22.200 91.600 26.200 ;
        RECT 96.000 22.200 96.800 27.800 ;
        RECT 100.400 27.400 101.000 30.400 ;
        RECT 105.600 28.400 106.200 31.800 ;
        RECT 106.800 28.800 107.600 30.400 ;
        RECT 103.600 27.600 106.200 28.400 ;
        RECT 108.400 28.200 109.200 28.400 ;
        RECT 107.600 27.600 109.200 28.200 ;
        RECT 98.800 26.800 101.000 27.400 ;
        RECT 98.800 22.200 99.600 26.800 ;
        RECT 103.800 26.200 104.400 27.600 ;
        RECT 107.600 27.200 108.400 27.600 ;
        RECT 105.400 26.200 109.000 26.600 ;
        RECT 103.600 22.200 104.400 26.200 ;
        RECT 105.200 26.000 109.200 26.200 ;
        RECT 105.200 22.200 106.000 26.000 ;
        RECT 108.400 22.200 109.200 26.000 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 6.000 15.000 6.800 19.800 ;
        RECT 10.400 18.400 11.200 19.800 ;
        RECT 9.200 17.800 11.200 18.400 ;
        RECT 14.800 17.800 15.600 19.800 ;
        RECT 19.000 18.400 20.200 19.800 ;
        RECT 18.800 17.800 20.200 18.400 ;
        RECT 9.200 17.000 10.000 17.800 ;
        RECT 14.800 17.200 15.400 17.800 ;
        RECT 12.600 16.600 15.400 17.200 ;
        RECT 18.800 17.000 19.600 17.800 ;
        RECT 12.600 16.400 13.400 16.600 ;
        RECT 20.600 15.400 21.400 15.600 ;
        RECT 23.600 15.400 24.400 19.800 ;
        RECT 25.200 15.800 26.000 19.800 ;
        RECT 26.800 16.000 27.600 19.800 ;
        RECT 30.000 16.000 30.800 19.800 ;
        RECT 38.000 16.300 38.800 19.800 ;
        RECT 26.800 15.800 30.800 16.000 ;
        RECT 20.600 14.800 24.400 15.400 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 4.400 11.600 5.200 13.200 ;
        RECT 18.800 12.800 19.600 13.000 ;
        RECT 8.200 12.400 9.000 12.600 ;
        RECT 8.200 11.800 13.200 12.400 ;
        RECT 18.800 12.200 22.600 12.800 ;
        RECT 21.800 12.000 22.600 12.200 ;
        RECT 12.400 11.600 13.200 11.800 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 20.200 11.400 21.000 11.600 ;
        RECT 23.600 11.400 24.400 14.800 ;
        RECT 25.400 14.400 26.000 15.800 ;
        RECT 27.000 15.400 30.600 15.800 ;
        RECT 31.700 15.700 38.800 16.300 ;
        RECT 29.200 14.400 30.000 14.800 ;
        RECT 25.200 13.600 27.800 14.400 ;
        RECT 29.200 14.300 30.800 14.400 ;
        RECT 31.700 14.300 32.300 15.700 ;
        RECT 29.200 13.800 32.300 14.300 ;
        RECT 30.000 13.700 32.300 13.800 ;
        RECT 30.000 13.600 30.800 13.700 ;
        RECT 27.200 12.400 27.800 13.600 ;
        RECT 26.800 11.600 27.800 12.400 ;
        RECT 28.400 11.600 29.200 13.200 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 6.000 11.000 11.600 11.200 ;
        RECT 6.000 10.800 11.800 11.000 ;
        RECT 20.200 10.800 24.400 11.400 ;
        RECT 6.000 10.600 15.800 10.800 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 6.000 2.200 6.800 10.600 ;
        RECT 11.000 10.200 15.800 10.600 ;
        RECT 9.200 9.000 14.600 9.600 ;
        RECT 9.200 8.800 10.000 9.000 ;
        RECT 13.800 8.800 14.600 9.000 ;
        RECT 15.200 9.000 15.800 10.200 ;
        RECT 16.600 9.000 17.400 9.200 ;
        RECT 15.200 8.400 17.400 9.000 ;
        RECT 12.600 7.400 13.400 7.600 ;
        RECT 15.400 7.400 16.200 7.600 ;
        RECT 9.200 6.200 10.000 7.000 ;
        RECT 12.600 6.800 16.200 7.400 ;
        RECT 14.800 6.200 15.400 6.800 ;
        RECT 18.800 6.200 19.600 7.000 ;
        RECT 9.200 5.600 11.200 6.200 ;
        RECT 10.400 2.200 11.200 5.600 ;
        RECT 14.800 2.200 15.600 6.200 ;
        RECT 19.000 2.200 20.200 6.200 ;
        RECT 23.600 2.200 24.400 10.800 ;
        RECT 25.200 10.200 26.000 10.400 ;
        RECT 27.200 10.200 27.800 11.600 ;
        RECT 25.200 9.600 26.600 10.200 ;
        RECT 27.200 9.600 28.200 10.200 ;
        RECT 26.000 8.400 26.600 9.600 ;
        RECT 26.000 7.600 26.800 8.400 ;
        RECT 27.400 2.200 28.200 9.600 ;
        RECT 38.000 2.200 38.800 15.700 ;
        RECT 39.600 15.600 40.400 17.200 ;
        RECT 41.800 16.400 42.600 19.800 ;
        RECT 41.800 15.800 43.600 16.400 ;
        RECT 39.600 10.300 40.400 10.400 ;
        RECT 41.200 10.300 42.000 10.400 ;
        RECT 39.600 9.700 42.000 10.300 ;
        RECT 39.600 9.600 40.400 9.700 ;
        RECT 41.200 8.800 42.000 9.700 ;
        RECT 42.800 10.300 43.600 15.800 ;
        RECT 47.200 14.400 48.000 19.800 ;
        RECT 55.000 16.400 56.600 19.800 ;
        RECT 54.000 15.800 56.600 16.400 ;
        RECT 60.400 15.800 61.200 19.800 ;
        RECT 62.000 16.000 62.800 19.800 ;
        RECT 65.200 16.000 66.000 19.800 ;
        RECT 62.000 15.800 66.000 16.000 ;
        RECT 67.400 16.400 68.200 19.800 ;
        RECT 67.400 15.800 69.200 16.400 ;
        RECT 54.000 15.600 56.200 15.800 ;
        RECT 47.200 14.200 48.400 14.400 ;
        RECT 46.200 13.600 48.400 14.200 ;
        RECT 54.000 13.600 54.800 14.400 ;
        RECT 46.200 10.400 46.800 13.600 ;
        RECT 54.200 13.200 54.800 13.600 ;
        RECT 54.200 12.400 55.000 13.200 ;
        RECT 55.600 12.400 56.200 15.600 ;
        RECT 60.600 14.400 61.200 15.800 ;
        RECT 62.200 15.400 65.800 15.800 ;
        RECT 57.200 14.300 58.000 14.400 ;
        RECT 60.400 14.300 63.000 14.400 ;
        RECT 57.200 13.700 63.000 14.300 ;
        RECT 57.200 12.800 58.000 13.700 ;
        RECT 60.400 13.600 63.000 13.700 ;
        RECT 48.400 11.600 50.000 12.400 ;
        RECT 44.400 10.300 45.200 10.400 ;
        RECT 42.800 9.700 45.200 10.300 ;
        RECT 42.800 2.200 43.600 9.700 ;
        RECT 44.400 9.600 45.200 9.700 ;
        RECT 46.000 9.600 46.800 10.400 ;
        RECT 50.800 9.600 51.600 11.200 ;
        RECT 52.400 10.800 53.200 12.400 ;
        RECT 55.600 11.600 56.400 12.400 ;
        RECT 58.800 12.300 59.600 12.400 ;
        RECT 60.400 12.300 61.200 12.400 ;
        RECT 58.800 12.200 61.200 12.300 ;
        RECT 58.000 11.700 61.200 12.200 ;
        RECT 58.000 11.600 59.600 11.700 ;
        RECT 60.400 11.600 61.200 11.700 ;
        RECT 55.600 11.400 56.200 11.600 ;
        RECT 54.200 10.800 56.200 11.400 ;
        RECT 58.000 11.200 58.800 11.600 ;
        RECT 54.200 10.200 54.800 10.800 ;
        RECT 60.400 10.200 61.200 10.400 ;
        RECT 62.400 10.200 63.000 13.600 ;
        RECT 63.600 12.300 64.400 13.200 ;
        RECT 63.600 11.700 67.500 12.300 ;
        RECT 63.600 11.600 64.400 11.700 ;
        RECT 66.900 10.400 67.500 11.700 ;
        RECT 46.200 7.000 46.800 9.600 ;
        RECT 47.600 7.600 48.400 9.200 ;
        RECT 46.200 6.400 49.800 7.000 ;
        RECT 46.200 6.200 46.800 6.400 ;
        RECT 46.000 2.200 46.800 6.200 ;
        RECT 49.200 6.200 49.800 6.400 ;
        RECT 49.200 2.200 50.000 6.200 ;
        RECT 52.400 2.800 53.200 10.200 ;
        RECT 54.000 3.400 54.800 10.200 ;
        RECT 55.600 9.600 59.600 10.200 ;
        RECT 60.400 9.600 61.800 10.200 ;
        RECT 62.400 9.600 63.400 10.200 ;
        RECT 55.600 2.800 56.400 9.600 ;
        RECT 52.400 2.200 56.400 2.800 ;
        RECT 58.800 2.200 59.600 9.600 ;
        RECT 61.200 8.400 61.800 9.600 ;
        RECT 61.200 7.600 62.000 8.400 ;
        RECT 62.600 2.200 63.400 9.600 ;
        RECT 66.800 8.800 67.600 10.400 ;
        RECT 68.400 2.200 69.200 15.800 ;
        RECT 70.000 10.300 70.800 10.400 ;
        RECT 71.600 10.300 72.400 19.800 ;
        RECT 81.200 15.000 82.000 19.800 ;
        RECT 85.600 18.400 86.400 19.800 ;
        RECT 84.400 17.800 86.400 18.400 ;
        RECT 90.000 17.800 90.800 19.800 ;
        RECT 94.200 18.400 95.400 19.800 ;
        RECT 94.000 17.800 95.400 18.400 ;
        RECT 84.400 17.000 85.200 17.800 ;
        RECT 90.000 17.200 90.600 17.800 ;
        RECT 87.800 16.600 90.600 17.200 ;
        RECT 94.000 17.000 94.800 17.800 ;
        RECT 87.800 16.400 88.600 16.600 ;
        RECT 95.800 15.400 96.600 15.600 ;
        RECT 98.800 15.400 99.600 19.800 ;
        RECT 95.800 14.800 99.600 15.400 ;
        RECT 94.000 12.800 94.800 13.000 ;
        RECT 83.400 12.400 84.200 12.600 ;
        RECT 83.400 11.800 88.400 12.400 ;
        RECT 94.000 12.200 97.800 12.800 ;
        RECT 97.000 12.000 97.800 12.200 ;
        RECT 98.800 12.300 99.600 14.800 ;
        RECT 100.400 15.200 101.200 19.800 ;
        RECT 106.800 18.300 107.600 19.800 ;
        RECT 108.400 18.300 109.200 18.400 ;
        RECT 106.800 17.700 109.200 18.300 ;
        RECT 105.200 15.600 106.000 17.200 ;
        RECT 100.400 14.600 102.600 15.200 ;
        RECT 100.400 12.300 101.200 13.200 ;
        RECT 87.600 11.600 88.400 11.800 ;
        RECT 98.800 11.700 101.200 12.300 ;
        RECT 95.400 11.400 96.200 11.600 ;
        RECT 98.800 11.400 99.600 11.700 ;
        RECT 100.400 11.600 101.200 11.700 ;
        RECT 102.000 11.600 102.600 14.600 ;
        RECT 70.000 9.700 72.400 10.300 ;
        RECT 70.000 9.600 70.800 9.700 ;
        RECT 71.600 2.200 72.400 9.700 ;
        RECT 81.200 11.000 86.800 11.200 ;
        RECT 81.200 10.800 87.000 11.000 ;
        RECT 95.400 10.800 99.600 11.400 ;
        RECT 81.200 10.600 91.000 10.800 ;
        RECT 81.200 2.200 82.000 10.600 ;
        RECT 86.200 10.200 91.000 10.600 ;
        RECT 84.400 9.000 89.800 9.600 ;
        RECT 84.400 8.800 85.200 9.000 ;
        RECT 89.000 8.800 89.800 9.000 ;
        RECT 90.400 9.000 91.000 10.200 ;
        RECT 91.800 9.000 92.600 9.200 ;
        RECT 90.400 8.400 92.600 9.000 ;
        RECT 87.800 7.400 88.600 7.600 ;
        RECT 90.600 7.400 91.400 7.600 ;
        RECT 84.400 6.200 85.200 7.000 ;
        RECT 87.800 6.800 91.400 7.400 ;
        RECT 90.000 6.200 90.600 6.800 ;
        RECT 94.000 6.200 94.800 7.000 ;
        RECT 84.400 5.600 86.400 6.200 ;
        RECT 85.600 2.200 86.400 5.600 ;
        RECT 90.000 2.200 90.800 6.200 ;
        RECT 94.200 2.200 95.400 6.200 ;
        RECT 98.800 2.200 99.600 10.800 ;
        RECT 102.000 10.800 103.200 11.600 ;
        RECT 102.000 10.200 102.600 10.800 ;
        RECT 100.400 9.600 102.600 10.200 ;
        RECT 100.400 2.200 101.200 9.600 ;
        RECT 106.800 2.200 107.600 17.700 ;
        RECT 108.400 17.600 109.200 17.700 ;
      LAYER metal2 ;
        RECT 1.200 66.200 2.000 71.800 ;
        RECT 4.400 64.200 5.200 75.800 ;
        RECT 7.600 69.600 8.400 70.400 ;
        RECT 14.000 64.200 14.800 75.800 ;
        RECT 38.000 69.600 38.800 70.400 ;
        RECT 44.400 69.600 45.200 70.400 ;
        RECT 49.200 69.600 50.000 70.400 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 18.800 65.600 19.600 66.400 ;
        RECT 30.000 65.600 30.800 66.400 ;
        RECT 18.900 64.400 19.500 65.600 ;
        RECT 18.800 63.600 19.600 64.400 ;
        RECT 20.400 63.600 21.200 64.400 ;
        RECT 1.200 50.200 2.000 55.800 ;
        RECT 4.400 46.200 5.200 57.800 ;
        RECT 7.600 51.600 8.400 52.400 ;
        RECT 7.700 44.400 8.300 51.600 ;
        RECT 14.000 46.200 14.800 57.800 ;
        RECT 18.800 57.600 19.600 58.400 ;
        RECT 17.200 51.600 18.000 52.400 ;
        RECT 4.400 43.600 5.200 44.400 ;
        RECT 7.600 43.600 8.400 44.400 ;
        RECT 4.500 38.400 5.100 43.600 ;
        RECT 7.600 39.600 8.400 40.400 ;
        RECT 2.800 37.600 3.600 38.400 ;
        RECT 4.400 37.600 5.200 38.400 ;
        RECT 2.900 34.400 3.500 37.600 ;
        RECT 2.800 33.600 3.600 34.400 ;
        RECT 6.000 33.600 6.800 34.400 ;
        RECT 6.100 32.400 6.700 33.600 ;
        RECT 7.700 32.400 8.300 39.600 ;
        RECT 17.300 34.400 17.900 51.600 ;
        RECT 20.500 46.400 21.100 63.600 ;
        RECT 38.100 58.400 38.700 69.600 ;
        RECT 42.800 65.600 43.600 66.400 ;
        RECT 55.600 65.600 56.400 66.400 ;
        RECT 42.900 58.400 43.500 65.600 ;
        RECT 50.800 63.600 51.600 64.400 ;
        RECT 58.800 63.600 59.600 64.400 ;
        RECT 63.600 63.600 64.400 64.400 ;
        RECT 50.900 58.400 51.500 63.600 ;
        RECT 38.000 57.600 38.800 58.400 ;
        RECT 42.800 57.600 43.600 58.400 ;
        RECT 50.800 57.600 51.600 58.400 ;
        RECT 41.200 55.600 42.000 56.400 ;
        RECT 41.300 54.400 41.900 55.600 ;
        RECT 42.900 54.400 43.500 57.600 ;
        RECT 46.000 55.600 46.800 56.400 ;
        RECT 46.100 54.400 46.700 55.600 ;
        RECT 25.200 53.600 26.000 54.400 ;
        RECT 34.800 53.600 35.600 54.400 ;
        RECT 36.400 53.600 37.200 54.400 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 42.800 53.600 43.600 54.400 ;
        RECT 46.000 53.600 46.800 54.400 ;
        RECT 22.000 51.600 22.800 52.400 ;
        RECT 23.600 51.600 24.400 52.400 ;
        RECT 22.100 50.400 22.700 51.600 ;
        RECT 22.000 49.600 22.800 50.400 ;
        RECT 20.400 45.600 21.200 46.400 ;
        RECT 20.500 40.400 21.100 45.600 ;
        RECT 20.400 39.600 21.200 40.400 ;
        RECT 22.100 38.400 22.700 49.600 ;
        RECT 23.700 38.400 24.300 51.600 ;
        RECT 25.300 50.400 25.900 53.600 ;
        RECT 34.900 50.400 35.500 53.600 ;
        RECT 36.500 52.400 37.100 53.600 ;
        RECT 36.400 51.600 37.200 52.400 ;
        RECT 44.400 51.600 45.200 52.400 ;
        RECT 25.200 49.600 26.000 50.400 ;
        RECT 33.200 49.600 34.000 50.400 ;
        RECT 34.800 49.600 35.600 50.400 ;
        RECT 22.000 37.600 22.800 38.400 ;
        RECT 23.600 37.600 24.400 38.400 ;
        RECT 20.400 35.600 21.200 36.400 ;
        RECT 41.200 35.600 42.000 36.400 ;
        RECT 14.000 33.600 14.800 34.400 ;
        RECT 17.200 33.600 18.000 34.400 ;
        RECT 20.500 32.400 21.100 35.600 ;
        RECT 41.300 34.400 41.900 35.600 ;
        RECT 26.800 33.600 27.600 34.400 ;
        RECT 30.000 33.600 30.800 34.400 ;
        RECT 41.200 33.600 42.000 34.400 ;
        RECT 6.000 31.600 6.800 32.400 ;
        RECT 7.600 31.600 8.400 32.400 ;
        RECT 14.000 31.600 14.800 32.400 ;
        RECT 20.400 31.600 21.200 32.400 ;
        RECT 25.200 31.600 26.000 32.400 ;
        RECT 25.300 30.400 25.900 31.600 ;
        RECT 4.400 29.600 5.200 30.400 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 25.200 29.600 26.000 30.400 ;
        RECT 26.900 28.400 27.500 33.600 ;
        RECT 14.000 27.600 14.800 28.400 ;
        RECT 26.800 27.600 27.600 28.400 ;
        RECT 14.100 26.400 14.700 27.600 ;
        RECT 30.100 26.400 30.700 33.600 ;
        RECT 44.500 32.400 45.100 51.600 ;
        RECT 47.600 49.600 48.400 50.400 ;
        RECT 47.600 47.600 48.400 48.400 ;
        RECT 47.700 38.400 48.300 47.600 ;
        RECT 47.600 37.600 48.400 38.400 ;
        RECT 50.900 34.400 51.500 57.600 ;
        RECT 57.200 53.600 58.000 54.400 ;
        RECT 58.900 52.400 59.500 63.600 ;
        RECT 63.700 56.400 64.300 63.600 ;
        RECT 63.600 55.600 64.400 56.400 ;
        RECT 60.400 53.600 61.200 54.400 ;
        RECT 58.800 51.600 59.600 52.400 ;
        RECT 52.400 45.600 53.200 46.400 ;
        RECT 52.500 34.400 53.100 45.600 ;
        RECT 54.000 43.600 54.800 44.400 ;
        RECT 54.100 38.400 54.700 43.600 ;
        RECT 54.000 37.600 54.800 38.400 ;
        RECT 50.800 33.600 51.600 34.400 ;
        RECT 52.400 33.600 53.200 34.400 ;
        RECT 44.400 31.600 45.200 32.400 ;
        RECT 46.000 27.600 46.800 28.400 ;
        RECT 14.000 25.600 14.800 26.400 ;
        RECT 23.600 25.600 24.400 26.400 ;
        RECT 30.000 25.600 30.800 26.400 ;
        RECT 23.700 24.400 24.300 25.600 ;
        RECT 23.600 23.600 24.400 24.400 ;
        RECT 28.400 23.600 29.200 24.400 ;
        RECT 41.200 23.600 42.000 24.400 ;
        RECT 49.200 23.600 50.000 24.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 4.500 10.400 5.100 11.600 ;
        RECT 4.400 9.600 5.200 10.400 ;
        RECT 6.000 10.200 6.800 15.800 ;
        RECT 9.200 6.200 10.000 17.800 ;
        RECT 12.400 11.600 13.200 12.400 ;
        RECT 18.800 6.200 19.600 17.800 ;
        RECT 25.200 15.600 26.000 16.400 ;
        RECT 25.300 10.400 25.900 15.600 ;
        RECT 28.500 12.400 29.100 23.600 ;
        RECT 39.600 15.600 40.400 16.400 ;
        RECT 26.800 11.600 27.600 12.400 ;
        RECT 28.400 11.600 29.200 12.400 ;
        RECT 39.700 10.400 40.300 15.600 ;
        RECT 23.600 9.600 24.400 10.400 ;
        RECT 25.200 9.600 26.000 10.400 ;
        RECT 39.600 9.600 40.400 10.400 ;
        RECT 23.700 8.400 24.300 9.600 ;
        RECT 41.300 8.400 41.900 23.600 ;
        RECT 47.600 13.600 48.400 14.400 ;
        RECT 49.300 12.400 49.900 23.600 ;
        RECT 52.500 12.400 53.100 33.600 ;
        RECT 60.500 32.400 61.100 53.600 ;
        RECT 65.300 36.400 65.900 69.600 ;
        RECT 66.800 65.600 67.600 66.400 ;
        RECT 78.000 66.200 78.800 71.800 ;
        RECT 66.900 54.400 67.500 65.600 ;
        RECT 81.200 64.200 82.000 75.800 ;
        RECT 84.400 69.600 85.200 70.400 ;
        RECT 73.200 55.600 74.000 56.400 ;
        RECT 66.800 53.600 67.600 54.400 ;
        RECT 68.400 53.600 69.200 54.400 ;
        RECT 68.500 52.400 69.100 53.600 ;
        RECT 68.400 51.600 69.200 52.400 ;
        RECT 70.000 51.600 70.800 52.400 ;
        RECT 71.600 49.600 72.400 50.400 ;
        RECT 73.300 48.400 73.900 55.600 ;
        RECT 76.400 53.600 77.200 54.400 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 78.000 51.600 78.800 52.400 ;
        RECT 78.100 50.400 78.700 51.600 ;
        RECT 78.000 49.600 78.800 50.400 ;
        RECT 81.200 49.600 82.000 50.400 ;
        RECT 73.200 47.600 74.000 48.400 ;
        RECT 81.300 38.400 81.900 49.600 ;
        RECT 84.500 38.400 85.100 69.600 ;
        RECT 90.800 64.200 91.600 75.800 ;
        RECT 98.800 71.800 99.600 72.600 ;
        RECT 105.400 71.800 106.200 72.600 ;
        RECT 98.800 68.400 99.400 71.800 ;
        RECT 102.800 68.400 103.600 68.600 ;
        RECT 98.800 67.800 103.600 68.400 ;
        RECT 98.800 67.000 99.400 67.800 ;
        RECT 105.600 67.000 106.200 71.800 ;
        RECT 98.800 66.200 99.600 67.000 ;
        RECT 105.400 66.200 106.200 67.000 ;
        RECT 95.600 63.600 96.400 64.400 ;
        RECT 100.400 63.600 101.200 64.400 ;
        RECT 94.000 57.600 94.800 58.400 ;
        RECT 94.100 56.400 94.700 57.600 ;
        RECT 89.200 55.600 90.000 56.400 ;
        RECT 94.000 55.600 94.800 56.400 ;
        RECT 95.600 55.600 96.400 56.400 ;
        RECT 100.500 56.300 101.100 63.600 ;
        RECT 98.900 55.700 101.100 56.300 ;
        RECT 89.300 54.400 89.900 55.600 ;
        RECT 89.200 53.600 90.000 54.400 ;
        RECT 89.300 52.400 89.900 53.600 ;
        RECT 89.200 51.600 90.000 52.400 ;
        RECT 94.100 48.400 94.700 55.600 ;
        RECT 95.700 52.400 96.300 55.600 ;
        RECT 97.200 53.600 98.000 54.400 ;
        RECT 95.600 51.600 96.400 52.400 ;
        RECT 94.000 47.600 94.800 48.400 ;
        RECT 94.000 43.600 94.800 44.400 ;
        RECT 81.200 37.600 82.000 38.400 ;
        RECT 84.400 37.600 85.200 38.400 ;
        RECT 65.200 35.600 66.000 36.400 ;
        RECT 76.400 35.600 77.200 36.400 ;
        RECT 60.400 31.600 61.200 32.400 ;
        RECT 54.000 29.600 54.800 30.400 ;
        RECT 54.100 28.400 54.700 29.600 ;
        RECT 54.000 27.600 54.800 28.400 ;
        RECT 57.200 27.600 58.000 28.400 ;
        RECT 54.000 15.600 54.800 16.400 ;
        RECT 54.000 13.600 54.800 14.400 ;
        RECT 60.500 12.400 61.100 31.600 ;
        RECT 65.300 30.400 65.900 35.600 ;
        RECT 94.100 34.400 94.700 43.600 ;
        RECT 98.900 36.400 99.500 55.700 ;
        RECT 100.400 53.600 101.200 54.400 ;
        RECT 100.500 48.400 101.100 53.600 ;
        RECT 102.000 51.600 102.800 52.400 ;
        RECT 105.200 51.600 106.000 52.400 ;
        RECT 105.300 50.400 105.900 51.600 ;
        RECT 103.600 49.600 104.400 50.400 ;
        RECT 105.200 49.600 106.000 50.400 ;
        RECT 100.400 47.600 101.200 48.400 ;
        RECT 102.000 47.600 102.800 48.400 ;
        RECT 100.400 45.600 101.200 46.400 ;
        RECT 102.100 42.300 102.700 47.600 ;
        RECT 103.700 44.400 104.300 49.600 ;
        RECT 105.200 47.600 106.000 48.400 ;
        RECT 106.800 47.600 107.600 48.400 ;
        RECT 105.300 46.400 105.900 47.600 ;
        RECT 106.900 46.400 107.500 47.600 ;
        RECT 105.200 45.600 106.000 46.400 ;
        RECT 106.800 45.600 107.600 46.400 ;
        RECT 103.600 43.600 104.400 44.400 ;
        RECT 100.500 41.700 102.700 42.300 ;
        RECT 95.600 35.600 96.400 36.400 ;
        RECT 98.800 35.600 99.600 36.400 ;
        RECT 95.700 34.400 96.300 35.600 ;
        RECT 73.200 33.600 74.000 34.400 ;
        RECT 92.400 33.600 93.200 34.400 ;
        RECT 94.000 33.600 94.800 34.400 ;
        RECT 95.600 33.600 96.400 34.400 ;
        RECT 73.300 32.400 73.900 33.600 ;
        RECT 92.500 32.400 93.100 33.600 ;
        RECT 95.700 32.400 96.300 33.600 ;
        RECT 70.000 31.600 70.800 32.400 ;
        RECT 73.200 31.600 74.000 32.400 ;
        RECT 92.400 31.600 93.200 32.400 ;
        RECT 95.600 31.600 96.400 32.400 ;
        RECT 97.200 31.600 98.000 32.400 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 71.600 29.600 72.400 30.400 ;
        RECT 87.600 29.600 88.400 30.400 ;
        RECT 94.000 29.600 94.800 30.400 ;
        RECT 98.800 29.600 99.600 30.400 ;
        RECT 71.700 28.400 72.300 29.600 ;
        RECT 68.400 27.600 69.200 28.400 ;
        RECT 71.600 27.600 72.400 28.400 ;
        RECT 87.700 26.400 88.300 29.600 ;
        RECT 94.100 28.400 94.700 29.600 ;
        RECT 90.800 27.600 91.600 28.400 ;
        RECT 94.000 27.600 94.800 28.400 ;
        RECT 84.400 25.600 85.200 26.400 ;
        RECT 87.600 25.600 88.400 26.400 ;
        RECT 84.500 20.400 85.100 25.600 ;
        RECT 84.400 19.600 85.200 20.400 ;
        RECT 98.800 19.600 99.600 20.400 ;
        RECT 98.900 18.400 99.500 19.600 ;
        RECT 49.200 11.600 50.000 12.400 ;
        RECT 52.400 11.600 53.200 12.400 ;
        RECT 60.400 11.600 61.200 12.400 ;
        RECT 68.400 11.600 69.200 12.400 ;
        RECT 44.400 9.600 45.200 10.400 ;
        RECT 50.800 9.600 51.600 10.400 ;
        RECT 60.400 9.600 61.200 10.400 ;
        RECT 66.800 9.600 67.600 10.400 ;
        RECT 70.000 9.600 70.800 10.400 ;
        RECT 81.200 10.200 82.000 15.800 ;
        RECT 23.600 7.600 24.400 8.400 ;
        RECT 41.200 7.600 42.000 8.400 ;
        RECT 47.600 7.600 48.400 8.400 ;
        RECT 84.400 6.200 85.200 17.800 ;
        RECT 87.600 11.600 88.400 12.400 ;
        RECT 94.000 6.200 94.800 17.800 ;
        RECT 98.800 17.600 99.600 18.400 ;
        RECT 100.500 12.400 101.100 41.700 ;
        RECT 105.200 41.600 106.000 42.400 ;
        RECT 103.600 31.600 104.400 32.400 ;
        RECT 105.300 30.400 105.900 41.600 ;
        RECT 106.800 37.600 107.600 38.400 ;
        RECT 106.800 33.600 107.600 34.400 ;
        RECT 106.900 30.400 107.500 33.600 ;
        RECT 105.200 29.600 106.000 30.400 ;
        RECT 106.800 29.600 107.600 30.400 ;
        RECT 105.300 16.400 105.900 29.600 ;
        RECT 108.400 27.600 109.200 28.400 ;
        RECT 108.500 26.400 109.100 27.600 ;
        RECT 108.400 25.600 109.200 26.400 ;
        RECT 108.500 18.400 109.100 25.600 ;
        RECT 108.400 17.600 109.200 18.400 ;
        RECT 105.200 15.600 106.000 16.400 ;
        RECT 100.400 11.600 101.200 12.400 ;
      LAYER metal3 ;
        RECT 7.600 70.300 8.400 70.400 ;
        RECT 38.000 70.300 38.800 70.400 ;
        RECT 7.600 69.700 38.800 70.300 ;
        RECT 7.600 69.600 8.400 69.700 ;
        RECT 38.000 69.600 38.800 69.700 ;
        RECT 44.400 70.300 45.200 70.400 ;
        RECT 49.200 70.300 50.000 70.400 ;
        RECT 44.400 69.700 50.000 70.300 ;
        RECT 44.400 69.600 45.200 69.700 ;
        RECT 49.200 69.600 50.000 69.700 ;
        RECT 18.800 66.300 19.600 66.400 ;
        RECT 30.000 66.300 30.800 66.400 ;
        RECT 55.600 66.300 56.400 66.400 ;
        RECT 66.800 66.300 67.600 66.400 ;
        RECT 18.800 65.700 67.600 66.300 ;
        RECT 18.800 65.600 19.600 65.700 ;
        RECT 30.000 65.600 30.800 65.700 ;
        RECT 55.600 65.600 56.400 65.700 ;
        RECT 66.800 65.600 67.600 65.700 ;
        RECT 95.600 64.300 96.400 64.400 ;
        RECT 100.400 64.300 101.200 64.400 ;
        RECT 95.600 63.700 101.200 64.300 ;
        RECT 95.600 63.600 96.400 63.700 ;
        RECT 100.400 63.600 101.200 63.700 ;
        RECT 18.800 58.300 19.600 58.400 ;
        RECT 42.800 58.300 43.600 58.400 ;
        RECT 18.800 57.700 43.600 58.300 ;
        RECT 18.800 57.600 19.600 57.700 ;
        RECT 42.800 57.600 43.600 57.700 ;
        RECT 50.800 58.300 51.600 58.400 ;
        RECT 94.000 58.300 94.800 58.400 ;
        RECT 50.800 57.700 94.800 58.300 ;
        RECT 50.800 57.600 51.600 57.700 ;
        RECT 94.000 57.600 94.800 57.700 ;
        RECT 41.200 56.300 42.000 56.400 ;
        RECT 46.000 56.300 46.800 56.400 ;
        RECT 41.200 55.700 46.800 56.300 ;
        RECT 41.200 55.600 42.000 55.700 ;
        RECT 46.000 55.600 46.800 55.700 ;
        RECT 63.600 56.300 64.400 56.400 ;
        RECT 89.200 56.300 90.000 56.400 ;
        RECT 95.600 56.300 96.400 56.400 ;
        RECT 63.600 55.700 88.300 56.300 ;
        RECT 63.600 55.600 64.400 55.700 ;
        RECT 25.200 54.300 26.000 54.400 ;
        RECT 34.800 54.300 35.600 54.400 ;
        RECT 25.200 53.700 35.600 54.300 ;
        RECT 25.200 53.600 26.000 53.700 ;
        RECT 34.800 53.600 35.600 53.700 ;
        RECT 42.800 54.300 43.600 54.400 ;
        RECT 57.200 54.300 58.000 54.400 ;
        RECT 68.400 54.300 69.200 54.400 ;
        RECT 76.400 54.300 77.200 54.400 ;
        RECT 42.800 53.700 77.200 54.300 ;
        RECT 87.700 54.300 88.300 55.700 ;
        RECT 89.200 55.700 96.400 56.300 ;
        RECT 89.200 55.600 90.000 55.700 ;
        RECT 95.600 55.600 96.400 55.700 ;
        RECT 97.200 54.300 98.000 54.400 ;
        RECT 87.700 53.700 98.000 54.300 ;
        RECT 42.800 53.600 43.600 53.700 ;
        RECT 57.200 53.600 58.000 53.700 ;
        RECT 68.400 53.600 69.200 53.700 ;
        RECT 76.400 53.600 77.200 53.700 ;
        RECT 97.200 53.600 98.000 53.700 ;
        RECT 17.200 52.300 18.000 52.400 ;
        RECT 36.400 52.300 37.200 52.400 ;
        RECT 70.000 52.300 70.800 52.400 ;
        RECT 17.200 51.700 70.800 52.300 ;
        RECT 17.200 51.600 18.000 51.700 ;
        RECT 36.400 51.600 37.200 51.700 ;
        RECT 70.000 51.600 70.800 51.700 ;
        RECT 74.800 52.300 75.600 52.400 ;
        RECT 89.200 52.300 90.000 52.400 ;
        RECT 74.800 51.700 90.000 52.300 ;
        RECT 74.800 51.600 75.600 51.700 ;
        RECT 89.200 51.600 90.000 51.700 ;
        RECT 94.000 52.300 94.800 52.400 ;
        RECT 102.000 52.300 102.800 52.400 ;
        RECT 94.000 51.700 102.800 52.300 ;
        RECT 94.000 51.600 94.800 51.700 ;
        RECT 102.000 51.600 102.800 51.700 ;
        RECT 22.000 50.300 22.800 50.400 ;
        RECT 33.200 50.300 34.000 50.400 ;
        RECT 22.000 49.700 34.000 50.300 ;
        RECT 22.000 49.600 22.800 49.700 ;
        RECT 33.200 49.600 34.000 49.700 ;
        RECT 34.800 50.300 35.600 50.400 ;
        RECT 47.600 50.300 48.400 50.400 ;
        RECT 34.800 49.700 48.400 50.300 ;
        RECT 34.800 49.600 35.600 49.700 ;
        RECT 47.600 49.600 48.400 49.700 ;
        RECT 71.600 50.300 72.400 50.400 ;
        RECT 78.000 50.300 78.800 50.400 ;
        RECT 71.600 49.700 78.800 50.300 ;
        RECT 71.600 49.600 72.400 49.700 ;
        RECT 78.000 49.600 78.800 49.700 ;
        RECT 81.200 50.300 82.000 50.400 ;
        RECT 105.200 50.300 106.000 50.400 ;
        RECT 81.200 49.700 106.000 50.300 ;
        RECT 81.200 49.600 82.000 49.700 ;
        RECT 105.200 49.600 106.000 49.700 ;
        RECT 47.600 48.300 48.400 48.400 ;
        RECT 73.200 48.300 74.000 48.400 ;
        RECT 47.600 47.700 74.000 48.300 ;
        RECT 47.600 47.600 48.400 47.700 ;
        RECT 73.200 47.600 74.000 47.700 ;
        RECT 94.000 48.300 94.800 48.400 ;
        RECT 100.400 48.300 101.200 48.400 ;
        RECT 94.000 47.700 101.200 48.300 ;
        RECT 94.000 47.600 94.800 47.700 ;
        RECT 100.400 47.600 101.200 47.700 ;
        RECT 102.000 48.300 102.800 48.400 ;
        RECT 105.200 48.300 106.000 48.400 ;
        RECT 102.000 47.700 106.000 48.300 ;
        RECT 102.000 47.600 102.800 47.700 ;
        RECT 105.200 47.600 106.000 47.700 ;
        RECT 20.400 46.300 21.200 46.400 ;
        RECT 52.400 46.300 53.200 46.400 ;
        RECT 20.400 45.700 53.200 46.300 ;
        RECT 20.400 45.600 21.200 45.700 ;
        RECT 52.400 45.600 53.200 45.700 ;
        RECT 100.400 46.300 101.200 46.400 ;
        RECT 106.800 46.300 107.600 46.400 ;
        RECT 100.400 45.700 107.600 46.300 ;
        RECT 100.400 45.600 101.200 45.700 ;
        RECT 106.800 45.600 107.600 45.700 ;
        RECT 4.400 44.300 5.200 44.400 ;
        RECT 7.600 44.300 8.400 44.400 ;
        RECT 4.400 43.700 8.400 44.300 ;
        RECT 4.400 43.600 5.200 43.700 ;
        RECT 7.600 43.600 8.400 43.700 ;
        RECT 54.000 44.300 54.800 44.400 ;
        RECT 103.600 44.300 104.400 44.400 ;
        RECT 54.000 43.700 104.400 44.300 ;
        RECT 54.000 43.600 54.800 43.700 ;
        RECT 103.600 43.600 104.400 43.700 ;
        RECT 100.400 42.300 101.200 42.400 ;
        RECT 105.200 42.300 106.000 42.400 ;
        RECT 100.400 41.700 106.000 42.300 ;
        RECT 100.400 41.600 101.200 41.700 ;
        RECT 105.200 41.600 106.000 41.700 ;
        RECT 7.600 40.300 8.400 40.400 ;
        RECT 20.400 40.300 21.200 40.400 ;
        RECT 7.600 39.700 21.200 40.300 ;
        RECT 7.600 39.600 8.400 39.700 ;
        RECT 20.400 39.600 21.200 39.700 ;
        RECT 2.800 38.300 3.600 38.400 ;
        RECT 23.600 38.300 24.400 38.400 ;
        RECT 2.800 37.700 24.400 38.300 ;
        RECT 2.800 37.600 3.600 37.700 ;
        RECT 23.600 37.600 24.400 37.700 ;
        RECT 84.400 38.300 85.200 38.400 ;
        RECT 106.800 38.300 107.600 38.400 ;
        RECT 84.400 37.700 107.600 38.300 ;
        RECT 84.400 37.600 85.200 37.700 ;
        RECT 106.800 37.600 107.600 37.700 ;
        RECT 20.400 36.300 21.200 36.400 ;
        RECT 41.200 36.300 42.000 36.400 ;
        RECT 20.400 35.700 42.000 36.300 ;
        RECT 20.400 35.600 21.200 35.700 ;
        RECT 41.200 35.600 42.000 35.700 ;
        RECT 65.200 36.300 66.000 36.400 ;
        RECT 76.400 36.300 77.200 36.400 ;
        RECT 65.200 35.700 77.200 36.300 ;
        RECT 65.200 35.600 66.000 35.700 ;
        RECT 76.400 35.600 77.200 35.700 ;
        RECT 95.600 36.300 96.400 36.400 ;
        RECT 98.800 36.300 99.600 36.400 ;
        RECT 95.600 35.700 99.600 36.300 ;
        RECT 95.600 35.600 96.400 35.700 ;
        RECT 98.800 35.600 99.600 35.700 ;
        RECT 6.000 34.300 6.800 34.400 ;
        RECT 14.000 34.300 14.800 34.400 ;
        RECT 6.000 33.700 14.800 34.300 ;
        RECT 6.000 33.600 6.800 33.700 ;
        RECT 14.000 33.600 14.800 33.700 ;
        RECT 17.200 34.300 18.000 34.400 ;
        RECT 26.800 34.300 27.600 34.400 ;
        RECT 17.200 33.700 27.600 34.300 ;
        RECT 17.200 33.600 18.000 33.700 ;
        RECT 26.800 33.600 27.600 33.700 ;
        RECT 30.000 34.300 30.800 34.400 ;
        RECT 50.800 34.300 51.600 34.400 ;
        RECT 30.000 33.700 51.600 34.300 ;
        RECT 30.000 33.600 30.800 33.700 ;
        RECT 50.800 33.600 51.600 33.700 ;
        RECT 52.400 34.300 53.200 34.400 ;
        RECT 92.400 34.300 93.200 34.400 ;
        RECT 52.400 33.700 93.200 34.300 ;
        RECT 52.400 33.600 53.200 33.700 ;
        RECT 92.400 33.600 93.200 33.700 ;
        RECT 94.000 34.300 94.800 34.400 ;
        RECT 106.800 34.300 107.600 34.400 ;
        RECT 94.000 33.700 107.600 34.300 ;
        RECT 94.000 33.600 94.800 33.700 ;
        RECT 106.800 33.600 107.600 33.700 ;
        RECT 14.000 32.300 14.800 32.400 ;
        RECT 25.200 32.300 26.000 32.400 ;
        RECT 44.400 32.300 45.200 32.400 ;
        RECT 14.000 31.700 45.200 32.300 ;
        RECT 14.000 31.600 14.800 31.700 ;
        RECT 25.200 31.600 26.000 31.700 ;
        RECT 44.400 31.600 45.200 31.700 ;
        RECT 60.400 32.300 61.200 32.400 ;
        RECT 70.000 32.300 70.800 32.400 ;
        RECT 60.400 31.700 70.800 32.300 ;
        RECT 60.400 31.600 61.200 31.700 ;
        RECT 70.000 31.600 70.800 31.700 ;
        RECT 73.200 32.300 74.000 32.400 ;
        RECT 95.600 32.300 96.400 32.400 ;
        RECT 73.200 31.700 96.400 32.300 ;
        RECT 73.200 31.600 74.000 31.700 ;
        RECT 95.600 31.600 96.400 31.700 ;
        RECT 97.200 32.300 98.000 32.400 ;
        RECT 103.600 32.300 104.400 32.400 ;
        RECT 97.200 31.700 104.400 32.300 ;
        RECT 97.200 31.600 98.000 31.700 ;
        RECT 103.600 31.600 104.400 31.700 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 7.600 30.300 8.400 30.400 ;
        RECT 4.400 29.700 8.400 30.300 ;
        RECT 4.400 29.600 5.200 29.700 ;
        RECT 7.600 29.600 8.400 29.700 ;
        RECT 98.800 30.300 99.600 30.400 ;
        RECT 105.200 30.300 106.000 30.400 ;
        RECT 98.800 29.700 106.000 30.300 ;
        RECT 98.800 29.600 99.600 29.700 ;
        RECT 105.200 29.600 106.000 29.700 ;
        RECT 14.000 28.300 14.800 28.400 ;
        RECT 46.000 28.300 46.800 28.400 ;
        RECT 14.000 27.700 46.800 28.300 ;
        RECT 14.000 27.600 14.800 27.700 ;
        RECT 46.000 27.600 46.800 27.700 ;
        RECT 54.000 28.300 54.800 28.400 ;
        RECT 57.200 28.300 58.000 28.400 ;
        RECT 54.000 27.700 58.000 28.300 ;
        RECT 54.000 27.600 54.800 27.700 ;
        RECT 57.200 27.600 58.000 27.700 ;
        RECT 68.400 28.300 69.200 28.400 ;
        RECT 71.600 28.300 72.400 28.400 ;
        RECT 68.400 27.700 72.400 28.300 ;
        RECT 68.400 27.600 69.200 27.700 ;
        RECT 71.600 27.600 72.400 27.700 ;
        RECT 90.800 28.300 91.600 28.400 ;
        RECT 94.000 28.300 94.800 28.400 ;
        RECT 90.800 27.700 94.800 28.300 ;
        RECT 90.800 27.600 91.600 27.700 ;
        RECT 94.000 27.600 94.800 27.700 ;
        RECT 87.600 26.300 88.400 26.400 ;
        RECT 108.400 26.300 109.200 26.400 ;
        RECT 87.600 25.700 109.200 26.300 ;
        RECT 87.600 25.600 88.400 25.700 ;
        RECT 108.400 25.600 109.200 25.700 ;
        RECT 23.600 24.300 24.400 24.400 ;
        RECT 49.200 24.300 50.000 24.400 ;
        RECT 23.600 23.700 50.000 24.300 ;
        RECT 23.600 23.600 24.400 23.700 ;
        RECT 49.200 23.600 50.000 23.700 ;
        RECT 84.400 20.300 85.200 20.400 ;
        RECT 94.000 20.300 94.800 20.400 ;
        RECT 98.800 20.300 99.600 20.400 ;
        RECT 84.400 19.700 99.600 20.300 ;
        RECT 84.400 19.600 85.200 19.700 ;
        RECT 94.000 19.600 94.800 19.700 ;
        RECT 98.800 19.600 99.600 19.700 ;
        RECT 25.200 16.300 26.000 16.400 ;
        RECT 54.000 16.300 54.800 16.400 ;
        RECT 25.200 15.700 54.800 16.300 ;
        RECT 25.200 15.600 26.000 15.700 ;
        RECT 54.000 15.600 54.800 15.700 ;
        RECT 47.600 14.300 48.400 14.400 ;
        RECT 54.000 14.300 54.800 14.400 ;
        RECT 47.600 13.700 54.800 14.300 ;
        RECT 47.600 13.600 48.400 13.700 ;
        RECT 54.000 13.600 54.800 13.700 ;
        RECT 12.400 12.300 13.200 12.400 ;
        RECT 26.800 12.300 27.600 12.400 ;
        RECT 12.400 11.700 27.600 12.300 ;
        RECT 12.400 11.600 13.200 11.700 ;
        RECT 26.800 11.600 27.600 11.700 ;
        RECT 49.200 12.300 50.000 12.400 ;
        RECT 68.400 12.300 69.200 12.400 ;
        RECT 49.200 11.700 69.200 12.300 ;
        RECT 49.200 11.600 50.000 11.700 ;
        RECT 68.400 11.600 69.200 11.700 ;
        RECT 87.600 12.300 88.400 12.400 ;
        RECT 100.400 12.300 101.200 12.400 ;
        RECT 87.600 11.700 101.200 12.300 ;
        RECT 87.600 11.600 88.400 11.700 ;
        RECT 100.400 11.600 101.200 11.700 ;
        RECT 4.400 10.300 5.200 10.400 ;
        RECT 23.600 10.300 24.400 10.400 ;
        RECT 39.600 10.300 40.400 10.400 ;
        RECT 4.400 9.700 40.400 10.300 ;
        RECT 4.400 9.600 5.200 9.700 ;
        RECT 23.600 9.600 24.400 9.700 ;
        RECT 39.600 9.600 40.400 9.700 ;
        RECT 44.400 10.300 45.200 10.400 ;
        RECT 50.800 10.300 51.600 10.400 ;
        RECT 60.400 10.300 61.200 10.400 ;
        RECT 44.400 9.700 61.200 10.300 ;
        RECT 44.400 9.600 45.200 9.700 ;
        RECT 50.800 9.600 51.600 9.700 ;
        RECT 60.400 9.600 61.200 9.700 ;
        RECT 66.800 10.300 67.600 10.400 ;
        RECT 70.000 10.300 70.800 10.400 ;
        RECT 66.800 9.700 70.800 10.300 ;
        RECT 66.800 9.600 67.600 9.700 ;
        RECT 70.000 9.600 70.800 9.700 ;
        RECT 41.200 8.300 42.000 8.400 ;
        RECT 47.600 8.300 48.400 8.400 ;
        RECT 41.200 7.700 48.400 8.300 ;
        RECT 41.200 7.600 42.000 7.700 ;
        RECT 47.600 7.600 48.400 7.700 ;
      LAYER metal4 ;
        RECT 93.800 19.400 95.000 52.600 ;
        RECT 100.200 41.400 101.400 64.600 ;
  END
END vending_machine_18105070
END LIBRARY

